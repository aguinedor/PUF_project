-- File generated automatically
-- Description : ROM including 256 random pairs
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity random_rom is
    Port (
        address : in  std_logic_vector(7 downto 0); -- Adresse sur 8 bits
        data_out : out std_logic_vector(15 downto 0) -- Données de sortie : 16 bits (2 x 8 bits)
    );
end random_rom;
architecture Behavioral of random_rom is
    type rom_type is array (0 to 255) of std_logic_vector(15 downto 0);
    constant ROM : rom_type := (
    0 => "01111000_01101001",
    1 => "00011100_11111011",
    2 => "10100101_01011010",
    3 => "11110111_11101101",
    4 => "01010010_01100010",
    5 => "00000101_11001010",
    6 => "01100110_11010011",
    7 => "00101111_11001100",
    8 => "10101011_01100101",
    9 => "00100111_00100101",
    10 => "00111001_00100011",
    11 => "01001000_10110010",
    12 => "00010101_11011100",
    13 => "11110101_01000000",
    14 => "10110100_11111101",
    15 => "10111000_01011100",
    16 => "00000011_11101000",
    17 => "10101000_00101110",
    18 => "11000001_10011101",
    19 => "01011010_00101100",
    20 => "11110001_00100010",
    21 => "11000010_11010101",
    22 => "11001011_00001100",
    23 => "10101100_00000100",
    24 => "10011011_10010011",
    25 => "00100100_11000001",
    26 => "01110101_10010001",
    27 => "10011001_10000110",
    28 => "00011010_01010010",
    29 => "11100111_10010111",
    30 => "00001100_00100110",
    31 => "00111011_11100100",
    32 => "10000110_11110111",
    33 => "10110110_11110000",
    34 => "01001011_00001110",
    35 => "11010011_11010110",
    36 => "01011111_01000011",
    37 => "01010001_10111111",
    38 => "01001110_10101110",
    39 => "11100010_11111000",
    40 => "10100110_10010101",
    41 => "10001000_01010110",
    42 => "11011101_10011001",
    43 => "00001110_01110000",
    44 => "10100111_11100111",
    45 => "11100110_11110100",
    46 => "10110101_01101100",
    47 => "01011110_01111000",
    48 => "10100011_00110101",
    49 => "01010110_10001110",
    50 => "01010101_00011111",
    51 => "11000101_11011111",
    52 => "11001010_00110110",
    53 => "11101010_11100101",
    54 => "10101010_00010010",
    55 => "10001110_11010010",
    56 => "01001001_01100100",
    57 => "01010000_01111001",
    58 => "10010111_01010001",
    59 => "00000001_01011011",
    60 => "10111101_00010000",
    61 => "01100100_10000001",
    62 => "00011001_00111010",
    63 => "11111101_00010111",
    64 => "01110100_00111111",
    65 => "00010010_10110001",
    66 => "11111001_10111100",
    67 => "00011110_11011000",
    68 => "01101100_11100001",
    69 => "00010001_10110111",
    70 => "10111010_11000110",
    71 => "01100000_00110111",
    72 => "00100001_10100000",
    73 => "10011010_10111000",
    74 => "11100100_00000101",
    75 => "01100011_01011110",
    76 => "01101011_11101100",
    77 => "00010100_01101010",
    78 => "01101111_11000101",
    79 => "10111100_01011101",
    80 => "10010110_00000000",
    81 => "00110100_01110001",
    82 => "00001000_00101011",
    83 => "11010110_11000111",
    84 => "00110000_00011110",
    85 => "11101011_01111111",
    86 => "00101010_11000011",
    87 => "00010110_00010001",
    88 => "00110110_11100011",
    89 => "10111110_01101101",
    90 => "10011101_00001000",
    91 => "10010101_11100000",
    92 => "00111100_00011101",
    93 => "01001101_01100000",
    94 => "00110111_11001101",
    95 => "10001101_00100001",
    96 => "01111001_01111011",
    97 => "01000100_10111101",
    98 => "01011001_00101111",
    99 => "11010100_10011111",
    100 => "10010010_00001111",
    101 => "01111010_01000010",
    102 => "00000110_10110110",
    103 => "11110110_00111110",
    104 => "10111001_10100001",
    105 => "01011101_00010011",
    106 => "11000011_01111110",
    107 => "10111111_01001110",
    108 => "00100011_00111101",
    109 => "10110001_11010100",
    110 => "11001111_11001111",
    111 => "11111011_01011111",
    112 => "10111011_00100100",
    113 => "01111100_10001101",
    114 => "01011100_10101011",
    115 => "00100000_00000011",
    116 => "10101101_11000010",
    117 => "11001100_11100010",
    118 => "01101001_01000101",
    119 => "00001101_11110110",
    120 => "10100000_01011001",
    121 => "11101110_01001010",
    122 => "10011111_11001001",
    123 => "11010000_00001011",
    124 => "10001111_10110100",
    125 => "01001111_10101001",
    126 => "10011100_11101011",
    127 => "11011011_10101010",
    128 => "10011110_11111111",
    129 => "00110011_10100100",
    130 => "10001001_00011011",
    131 => "10010000_11000000",
    132 => "11000100_01010100",
    133 => "01100101_10000000",
    134 => "11110011_01110011",
    135 => "00010000_10011110",
    136 => "00000000_10101111",
    137 => "10010100_00110100",
    138 => "11010001_10010000",
    139 => "01011011_01010000",
    140 => "11101000_10111001",
    141 => "01111011_11011011",
    142 => "01110001_00110010",
    143 => "11000110_01100001",
    144 => "10000010_10100010",
    145 => "00111000_10011100",
    146 => "00101101_00010101",
    147 => "10001010_00011001",
    148 => "11111010_00000111",
    149 => "00011000_10001010",
    150 => "11011001_10000010",
    151 => "10110010_00010100",
    152 => "11101100_11101111",
    153 => "11111100_01001101",
    154 => "11110010_10110011",
    155 => "00010011_01001000",
    156 => "00101100_10100011",
    157 => "00101011_00101001",
    158 => "00000010_01101000",
    159 => "10001011_10010110",
    160 => "11001110_01101111",
    161 => "01101110_00010110",
    162 => "01110010_10101100",
    163 => "10101111_11101110",
    164 => "00100110_10001111",
    165 => "01001010_00100111",
    166 => "00011011_10000011",
    167 => "10011000_11111100",
    168 => "10000101_00101101",
    169 => "00101000_00001101",
    170 => "10100100_11010001",
    171 => "11010101_00111000",
    172 => "11111110_10111010",
    173 => "01101000_10100111",
    174 => "01101101_11101010",
    175 => "10110000_00011100",
    176 => "00110001_10101101",
    177 => "11110100_01000110",
    178 => "00110010_10011000",
    179 => "11011010_01110111",
    180 => "01010100_10001011",
    181 => "01000110_01110010",
    182 => "00000111_00110011",
    183 => "11111111_00111100",
    184 => "11001101_10001000",
    185 => "00100101_11011001",
    186 => "11000111_00111001",
    187 => "11101111_10011010",
    188 => "11001001_11111010",
    189 => "00111010_00000110",
    190 => "01111111_00000001",
    191 => "01011000_11011010",
    192 => "01110000_01011000",
    193 => "11010111_00000010",
    194 => "00111101_11000100",
    195 => "11111000_01000001",
    196 => "11110000_11010111",
    197 => "11011100_11111110",
    198 => "10101110_10110000",
    199 => "00111111_10110101",
    200 => "01000000_01100111",
    201 => "00000100_00001010",
    202 => "01000011_00101010",
    203 => "11011111_01010111",
    204 => "01001100_01001011",
    205 => "01111110_11011110",
    206 => "11100101_10001100",
    207 => "01110110_00001001",
    208 => "10001100_00100000",
    209 => "10000001_11001000",
    210 => "01100111_10010100",
    211 => "00001010_11001110",
    212 => "00001011_11111001",
    213 => "01101010_01010011",
    214 => "11011000_01001100",
    215 => "00010111_10100110",
    216 => "01000010_00011000",
    217 => "10101001_10100101",
    218 => "00101110_10010010",
    219 => "00001111_11010000",
    220 => "00100010_01100011",
    221 => "10000000_11001011",
    222 => "01000001_00111011",
    223 => "01010111_01110101",
    224 => "11011110_11110011",
    225 => "10100010_00110001",
    226 => "00111110_00101000",
    227 => "10000100_11100110",
    228 => "01111101_01101110",
    229 => "01000101_01001001",
    230 => "00110101_11011101",
    231 => "01010011_00110000",
    232 => "00101001_11110101",
    233 => "01110111_10001001",
    234 => "01100001_11110001",
    235 => "11100011_01111100",
    236 => "10000111_10101000",
    237 => "10010011_01010101",
    238 => "01000111_01110110",
    239 => "11101101_10000100",
    240 => "11100001_00011010",
    241 => "11000000_10111110",
    242 => "10100001_10111011",
    243 => "10110111_01100110",
    244 => "10010001_01111101",
    245 => "11101001_10011011",
    246 => "11001000_11110010",
    247 => "11100000_10000101",
    248 => "01100010_10000111",
    249 => "00001001_01111010",
    250 => "10110011_01101011",
    251 => "01110011_01001111",
    252 => "00011101_01110100",
    253 => "11010010_11101001",
    254 => "10000011_01000111",
    255 => "00011111_01000100"
    others => (others => '0')
    );
begin
    process(address)
    begin
        if (to_integer(unsigned(address)) <= 255) then
            data_out <= ROM(to_integer(unsigned(address)));
        else
            data_out <= (others => '0');
        end if;
    end process;
end Behavioral;
