-- File generated automatically
-- Description : ROM including 256 random pairs
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity random_rom is
    Port (
        address : integer range 0 to 255; -- Adresse sur 8 bits
        data_out : out std_logic_vector(15 downto 0) -- Données de sortie : 16 bits (2 x 8 bits)
    );
end random_rom;
architecture Behavioral of random_rom is
    type rom_type is array (0 to 255) of std_logic_vector(15 downto 0);
    constant ROM : rom_type := (
    0 => "0001001000000101",
    1 => "1100110000101111",
    2 => "1000110100111101",
    3 => "0110001101010010",
    4 => "1110101010110010",
    5 => "1011101001100010",
    6 => "0010011011100101",
    7 => "0000101010001101",
    8 => "0010101101001000",
    9 => "1001111111001010",
    10 => "0010110011010010",
    11 => "0001100110001111",
    12 => "1110110111000011",
    13 => "1100100101101011",
    14 => "0111110010000101",
    15 => "0000111101101101",
    16 => "0010100111101111",
    17 => "0100001001011011",
    18 => "1001101100001011",
    19 => "0101101111110010",
    20 => "1011110000110100",
    21 => "1100100001110000",
    22 => "0000001000011100",
    23 => "1000011011010011",
    24 => "0011101110110000",
    25 => "1100101011010001",
    26 => "1111100011010101",
    27 => "0111100110010001",
    28 => "1111001111001110",
    29 => "0000110101010110",
    30 => "1101010010101101",
    31 => "0110100110010100",
    32 => "1001001101100101",
    33 => "1111100100011110",
    34 => "1101001010101111",
    35 => "0101001001010001",
    36 => "0001101001001110",
    37 => "1110101101001100",
    38 => "1100111101001111",
    39 => "0010101010011101",
    40 => "1011001011000010",
    41 => "0101000001011101",
    42 => "0100101101100000",
    43 => "1000000111110011",
    44 => "0000000010110110",
    45 => "1001100001010111",
    46 => "0011000100100101",
    47 => "0001001100010001",
    48 => "0101101011011101",
    49 => "1100001100011011",
    50 => "1001111010100111",
    51 => "1101111110011011",
    52 => "1111010001000110",
    53 => "1101101111010100",
    54 => "0010111001110001",
    55 => "1001110100111000",
    56 => "1000101000110000",
    57 => "1010100101000010",
    58 => "0011011011010111",
    59 => "0011101010010011",
    60 => "1010101010111100",
    61 => "1010001101010101",
    62 => "0000011010000011",
    63 => "1110011101110011",
    64 => "1111011110011110",
    65 => "0011011110011111",
    66 => "0001101100101000",
    67 => "1000001100010110",
    68 => "0100011110110100",
    69 => "0000111011100100",
    70 => "1000110010000110",
    71 => "0110000011111100",
    72 => "1101111010101011",
    73 => "1010000000010011",
    74 => "0000100011110110",
    75 => "0011111000010010",
    76 => "1011100010101010",
    77 => "1101110100010111",
    78 => "1000001011101110",
    79 => "1110110010010111",
    80 => "0011010011111101",
    81 => "1000100010010110",
    82 => "1010011000110111",
    83 => "0110001000101101",
    84 => "1011011110111000",
    85 => "1100000101100111",
    86 => "1100101100011010",
    87 => "0100010111101001",
    88 => "0011110111110001",
    89 => "1100011000101110",
    90 => "1100011100001100",
    91 => "0110110111101101",
    92 => "1010111010011100",
    93 => "1001100111100010",
    94 => "1010011111111001",
    95 => "0100000000101001",
    96 => "1011101110001100",
    97 => "0001110111101000",
    98 => "0110101010001000",
    99 => "0011010110100010",
    100 => "0100001111111011",
    101 => "1010111100100001",
    102 => "0010111101001101",
    103 => "0000101100100110",
    104 => "0111011101001010",
    105 => "1101010100010100",
    106 => "0111010100000111",
    107 => "0001000110111010",
    108 => "0100110111000001",
    109 => "1111000101101000",
    110 => "0100000100000110",
    111 => "1111010111011011",
    112 => "0100111100101011",
    113 => "1100010111001001",
    114 => "0001010101111011",
    115 => "1011010100111100",
    116 => "0100111010000010",
    117 => "1011100101111100",
    118 => "0111110111111110",
    119 => "1011010001000011",
    120 => "1001010001011010",
    121 => "0111100001000100",
    122 => "0110111011101100",
    123 => "1010101110000000",
    124 => "1111000011011110",
    125 => "1100110100001000",
    126 => "0010000011110101",
    127 => "0001100011001101",
    128 => "0101111000000000",
    129 => "0100101011110000",
    130 => "1110100100000100",
    131 => "1101011000100000",
    132 => "1011011010101001",
    133 => "1000000000110010",
    134 => "0111101100110101",
    135 => "0001111111000100",
    136 => "1001001010100001",
    137 => "0001011111111010",
    138 => "0100010001000000",
    139 => "0101010111001011",
    140 => "0101000110111111",
    141 => "1011111000001110",
    142 => "1001000110011010",
    143 => "0010110110110011",
    144 => "1110000011111111",
    145 => "1010000111100111",
    146 => "0110101110011001",
    147 => "1111011000101100",
    148 => "0101011001101001",
    149 => "1110000110001001",
    150 => "0101010011001000",
    151 => "1000011101000101",
    152 => "1100111011001100",
    153 => "0001111001011001",
    154 => "0010010001100011",
    155 => "0111111101110100",
    156 => "0000011101011111",
    157 => "1101001110100000",
    158 => "1101110011011001",
    159 => "0011100001001001",
    160 => "1011001101101100",
    161 => "1000010001100001",
    162 => "0000100101111010",
    163 => "0010100000000011",
    164 => "1010010110100110",
    165 => "1111111101110010",
    166 => "1110001101001011",
    167 => "1101000010101110",
    168 => "1010110100110001",
    169 => "0000000101010000",
    170 => "0111000001111110",
    171 => "1111110101110101",
    172 => "0100110000011000",
    173 => "1000100110101000",
    174 => "1010001000101010",
    175 => "0110011011011100",
    176 => "1110111010110001",
    177 => "0111011010100100",
    178 => "0100011001111101",
    179 => "0001011010000111",
    180 => "1111101110001011",
    181 => "1110010111101011",
    182 => "1011110111000000",
    183 => "1111110010100011",
    184 => "1000101100100100",
    185 => "1110111110111101",
    186 => "1110011001000001",
    187 => "0011001100010000",
    188 => "1110100000111010",
    189 => "1001011111001111",
    190 => "0111101010111001",
    191 => "0101100111110100",
    192 => "1010110001101110",
    193 => "1011000100001010",
    194 => "0101110010000001",
    195 => "0011111111100001",
    196 => "0101001101100100",
    197 => "1101100100001111",
    198 => "1010100000000010",
    199 => "0110110001010100",
    200 => "0111001000111011",
    201 => "1001110001011100",
    202 => "0001010000011001",
    203 => "1001011001101111",
    204 => "1111101000111110",
    205 => "1001010111101010",
    206 => "0000110010110101",
    207 => "1000010100111111",
    208 => "0111001101110111",
    209 => "0001110001000111",
    210 => "1000111101111111",
    211 => "0010000111010000",
    212 => "0111000101101010",
    213 => "0010010110000100",
    214 => "0111111000001101",
    215 => "0100100110010101",
    216 => "1100001000100011",
    217 => "1001000000100010",
    218 => "0011000001110110",
    219 => "0100100001100110",
    220 => "0101111110001010",
    221 => "1100000000011101",
    222 => "0000010110101100",
    223 => "0110000101011000",
    224 => "1100010000110011",
    225 => "0110111110001110",
    226 => "0011100100110110",
    227 => "0000001111000111",
    228 => "1110010001111001",
    229 => "1000111011110111",
    230 => "0111010011011010",
    231 => "1111111001111000",
    232 => "1101100000000001",
    233 => "1011111101011110",
    234 => "1001101011011000",
    235 => "0110100010110111",
    236 => "0010001010111011",
    237 => "1101011110010010",
    238 => "0110010011000110",
    239 => "0011110010011000",
    240 => "1110001000011111",
    241 => "1101101010010000",
    242 => "1010010000100111",
    243 => "1101000110111110",
    244 => "0000010000001001",
    245 => "0110010101010011",
    246 => "0101011100111001",
    247 => "0001000010100101",
    248 => "0110011111011111",
    249 => "0101100011010110",
    250 => "1111001011100000",
    251 => "0011001000010101",
    252 => "0101110111100110",
    253 => "0010011111111000",
    254 => "0010001111000101",
    255 => "1011000011100011"
    );
begin
    process(address)
    begin
        data_out <= ROM(address);
    end process;
end Behavioral;
