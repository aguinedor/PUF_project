module ring_oscillator
  (input  enable,
   output ro_out);
  reg [6:0] inverters;
  (* KEEP="TRUE" *) wire nand_out;
  (* KEEP="TRUE" *) wire n11036_o;
  (* KEEP="TRUE" *) wire n11037_o;
  (* KEEP="TRUE" *) wire n11042_o;
  (* KEEP="TRUE" *) wire n11046_o;
  (* KEEP="TRUE" *) wire n11049_o;
  (* KEEP="TRUE" *) wire n11053_o;
  (* KEEP="TRUE" *) wire n11056_o;
  (* KEEP="TRUE" *) wire n11060_o;
  (* KEEP="TRUE" *) wire n11063_o;
  (* KEEP="TRUE" *) wire n11067_o;
  (* KEEP="TRUE" *) wire n11070_o;
  (* KEEP="TRUE" *) wire n11074_o;
  (* KEEP="TRUE" *) wire n11077_o;
  (* KEEP="TRUE" *) wire n11081_o;
  (* KEEP="TRUE" *) wire n11084_o;
  (* KEEP="TRUE" *) wire n11086_o;
  (* KEEP="TRUE" *) wire [6:0] n11087_o;
  assign ro_out = n11086_o;
  /* RTL_PUF/vhdl/ring_oscillator_no_lut.vhd:16:12  */
  always @*
    inverters = n11087_o; // (isignal)
  initial
    inverters = 7'b0000000;
  /* RTL_PUF/vhdl/ring_oscillator_no_lut.vhd:17:12  */
  assign nand_out = n11037_o; // (signal)
  /* RTL_PUF/vhdl/ring_oscillator_no_lut.vhd:24:38  */
  assign n11036_o = inverters[5];
  /* RTL_PUF/vhdl/ring_oscillator_no_lut.vhd:24:24  */
  assign n11037_o = ~(enable & n11036_o);
  /* RTL_PUF/vhdl/ring_oscillator_no_lut.vhd:29:9  */
  assign n11042_o = nand_out ? 1'b0 : 1'b1;
  /* RTL_PUF/vhdl/ring_oscillator_no_lut.vhd:40:25  */
  assign n11046_o = inverters[0];
  /* RTL_PUF/vhdl/ring_oscillator_no_lut.vhd:40:13  */
  assign n11049_o = n11046_o ? 1'b0 : 1'b1;
  /* RTL_PUF/vhdl/ring_oscillator_no_lut.vhd:40:25  */
  assign n11053_o = inverters[1];
  /* RTL_PUF/vhdl/ring_oscillator_no_lut.vhd:40:13  */
  assign n11056_o = n11053_o ? 1'b0 : 1'b1;
  /* RTL_PUF/vhdl/ring_oscillator_no_lut.vhd:40:25  */
  assign n11060_o = inverters[2];
  /* RTL_PUF/vhdl/ring_oscillator_no_lut.vhd:40:13  */
  assign n11063_o = n11060_o ? 1'b0 : 1'b1;
  /* RTL_PUF/vhdl/ring_oscillator_no_lut.vhd:40:25  */
  assign n11067_o = inverters[3];
  /* RTL_PUF/vhdl/ring_oscillator_no_lut.vhd:40:13  */
  assign n11070_o = n11067_o ? 1'b0 : 1'b1;
  /* RTL_PUF/vhdl/ring_oscillator_no_lut.vhd:40:25  */
  assign n11074_o = inverters[4];
  /* RTL_PUF/vhdl/ring_oscillator_no_lut.vhd:40:13  */
  assign n11077_o = n11074_o ? 1'b0 : 1'b1;
  /* RTL_PUF/vhdl/ring_oscillator_no_lut.vhd:40:25  */
  assign n11081_o = inverters[5];
  /* RTL_PUF/vhdl/ring_oscillator_no_lut.vhd:40:13  */
  assign n11084_o = n11081_o ? 1'b0 : 1'b1;
  /* RTL_PUF/vhdl/ring_oscillator_no_lut.vhd:49:24  */
  assign n11086_o = inverters[6];
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  assign n11087_o = {n11084_o, n11077_o, n11070_o, n11063_o, n11056_o, n11049_o, n11042_o};
endmodule

module random_rom
  (input  [7:0] address,
   output [15:0] data_out);
  (* KEEP="TRUE" *) wire [7:0] n11027_o;
  (* KEEP="TRUE" *) wire [15:0] n11033_data; // mem_rd
  assign data_out = n11033_data;
  /* RTL_PUF/vhdl/random_rom.vhd:275:25  */
  assign n11027_o = 8'b11111111 - address;
  /* RTL_PUF/vhdl/random_rom.vhd:9:9  */
  (* KEEP="TRUE" *) reg [15:0] n11032[255:0] ; // memory
  initial begin
    n11032[255] = 16'b0001001000000101;
    n11032[254] = 16'b1100110000101111;
    n11032[253] = 16'b1000110100111101;
    n11032[252] = 16'b0110001101010010;
    n11032[251] = 16'b1110101010110010;
    n11032[250] = 16'b1011101001100010;
    n11032[249] = 16'b0010011011100101;
    n11032[248] = 16'b0000101010001101;
    n11032[247] = 16'b0010101101001000;
    n11032[246] = 16'b1001111111001010;
    n11032[245] = 16'b0010110011010010;
    n11032[244] = 16'b0001100110001111;
    n11032[243] = 16'b1110110111000011;
    n11032[242] = 16'b1100100101101011;
    n11032[241] = 16'b0111110010000101;
    n11032[240] = 16'b0000111101101101;
    n11032[239] = 16'b0010100111101111;
    n11032[238] = 16'b0100001001011011;
    n11032[237] = 16'b1001101100001011;
    n11032[236] = 16'b0101101111110010;
    n11032[235] = 16'b1011110000110100;
    n11032[234] = 16'b1100100001110000;
    n11032[233] = 16'b0000001000011100;
    n11032[232] = 16'b1000011011010011;
    n11032[231] = 16'b0011101110110000;
    n11032[230] = 16'b1100101011010001;
    n11032[229] = 16'b1111100011010101;
    n11032[228] = 16'b0111100110010001;
    n11032[227] = 16'b1111001111001110;
    n11032[226] = 16'b0000110101010110;
    n11032[225] = 16'b1101010010101101;
    n11032[224] = 16'b0110100110010100;
    n11032[223] = 16'b1001001101100101;
    n11032[222] = 16'b1111100100011110;
    n11032[221] = 16'b1101001010101111;
    n11032[220] = 16'b0101001001010001;
    n11032[219] = 16'b0001101001001110;
    n11032[218] = 16'b1110101101001100;
    n11032[217] = 16'b1100111101001111;
    n11032[216] = 16'b0010101010011101;
    n11032[215] = 16'b1011001011000010;
    n11032[214] = 16'b0101000001011101;
    n11032[213] = 16'b0100101101100000;
    n11032[212] = 16'b1000000111110011;
    n11032[211] = 16'b0000000010110110;
    n11032[210] = 16'b1001100001010111;
    n11032[209] = 16'b0011000100100101;
    n11032[208] = 16'b0001001100010001;
    n11032[207] = 16'b0101101011011101;
    n11032[206] = 16'b1100001100011011;
    n11032[205] = 16'b1001111010100111;
    n11032[204] = 16'b1101111110011011;
    n11032[203] = 16'b1111010001000110;
    n11032[202] = 16'b1101101111010100;
    n11032[201] = 16'b0010111001110001;
    n11032[200] = 16'b1001110100111000;
    n11032[199] = 16'b1000101000110000;
    n11032[198] = 16'b1010100101000010;
    n11032[197] = 16'b0011011011010111;
    n11032[196] = 16'b0011101010010011;
    n11032[195] = 16'b1010101010111100;
    n11032[194] = 16'b1010001101010101;
    n11032[193] = 16'b0000011010000011;
    n11032[192] = 16'b1110011101110011;
    n11032[191] = 16'b1111011110011110;
    n11032[190] = 16'b0011011110011111;
    n11032[189] = 16'b0001101100101000;
    n11032[188] = 16'b1000001100010110;
    n11032[187] = 16'b0100011110110100;
    n11032[186] = 16'b0000111011100100;
    n11032[185] = 16'b1000110010000110;
    n11032[184] = 16'b0110000011111100;
    n11032[183] = 16'b1101111010101011;
    n11032[182] = 16'b1010000000010011;
    n11032[181] = 16'b0000100011110110;
    n11032[180] = 16'b0011111000010010;
    n11032[179] = 16'b1011100010101010;
    n11032[178] = 16'b1101110100010111;
    n11032[177] = 16'b1000001011101110;
    n11032[176] = 16'b1110110010010111;
    n11032[175] = 16'b0011010011111101;
    n11032[174] = 16'b1000100010010110;
    n11032[173] = 16'b1010011000110111;
    n11032[172] = 16'b0110001000101101;
    n11032[171] = 16'b1011011110111000;
    n11032[170] = 16'b1100000101100111;
    n11032[169] = 16'b1100101100011010;
    n11032[168] = 16'b0100010111101001;
    n11032[167] = 16'b0011110111110001;
    n11032[166] = 16'b1100011000101110;
    n11032[165] = 16'b1100011100001100;
    n11032[164] = 16'b0110110111101101;
    n11032[163] = 16'b1010111010011100;
    n11032[162] = 16'b1001100111100010;
    n11032[161] = 16'b1010011111111001;
    n11032[160] = 16'b0100000000101001;
    n11032[159] = 16'b1011101110001100;
    n11032[158] = 16'b0001110111101000;
    n11032[157] = 16'b0110101010001000;
    n11032[156] = 16'b0011010110100010;
    n11032[155] = 16'b0100001111111011;
    n11032[154] = 16'b1010111100100001;
    n11032[153] = 16'b0010111101001101;
    n11032[152] = 16'b0000101100100110;
    n11032[151] = 16'b0111011101001010;
    n11032[150] = 16'b1101010100010100;
    n11032[149] = 16'b0111010100000111;
    n11032[148] = 16'b0001000110111010;
    n11032[147] = 16'b0100110111000001;
    n11032[146] = 16'b1111000101101000;
    n11032[145] = 16'b0100000100000110;
    n11032[144] = 16'b1111010111011011;
    n11032[143] = 16'b0100111100101011;
    n11032[142] = 16'b1100010111001001;
    n11032[141] = 16'b0001010101111011;
    n11032[140] = 16'b1011010100111100;
    n11032[139] = 16'b0100111010000010;
    n11032[138] = 16'b1011100101111100;
    n11032[137] = 16'b0111110111111110;
    n11032[136] = 16'b1011010001000011;
    n11032[135] = 16'b1001010001011010;
    n11032[134] = 16'b0111100001000100;
    n11032[133] = 16'b0110111011101100;
    n11032[132] = 16'b1010101110000000;
    n11032[131] = 16'b1111000011011110;
    n11032[130] = 16'b1100110100001000;
    n11032[129] = 16'b0010000011110101;
    n11032[128] = 16'b0001100011001101;
    n11032[127] = 16'b0101111000000000;
    n11032[126] = 16'b0100101011110000;
    n11032[125] = 16'b1110100100000100;
    n11032[124] = 16'b1101011000100000;
    n11032[123] = 16'b1011011010101001;
    n11032[122] = 16'b1000000000110010;
    n11032[121] = 16'b0111101100110101;
    n11032[120] = 16'b0001111111000100;
    n11032[119] = 16'b1001001010100001;
    n11032[118] = 16'b0001011111111010;
    n11032[117] = 16'b0100010001000000;
    n11032[116] = 16'b0101010111001011;
    n11032[115] = 16'b0101000110111111;
    n11032[114] = 16'b1011111000001110;
    n11032[113] = 16'b1001000110011010;
    n11032[112] = 16'b0010110110110011;
    n11032[111] = 16'b1110000011111111;
    n11032[110] = 16'b1010000111100111;
    n11032[109] = 16'b0110101110011001;
    n11032[108] = 16'b1111011000101100;
    n11032[107] = 16'b0101011001101001;
    n11032[106] = 16'b1110000110001001;
    n11032[105] = 16'b0101010011001000;
    n11032[104] = 16'b1000011101000101;
    n11032[103] = 16'b1100111011001100;
    n11032[102] = 16'b0001111001011001;
    n11032[101] = 16'b0010010001100011;
    n11032[100] = 16'b0111111101110100;
    n11032[99] = 16'b0000011101011111;
    n11032[98] = 16'b1101001110100000;
    n11032[97] = 16'b1101110011011001;
    n11032[96] = 16'b0011100001001001;
    n11032[95] = 16'b1011001101101100;
    n11032[94] = 16'b1000010001100001;
    n11032[93] = 16'b0000100101111010;
    n11032[92] = 16'b0010100000000011;
    n11032[91] = 16'b1010010110100110;
    n11032[90] = 16'b1111111101110010;
    n11032[89] = 16'b1110001101001011;
    n11032[88] = 16'b1101000010101110;
    n11032[87] = 16'b1010110100110001;
    n11032[86] = 16'b0000000101010000;
    n11032[85] = 16'b0111000001111110;
    n11032[84] = 16'b1111110101110101;
    n11032[83] = 16'b0100110000011000;
    n11032[82] = 16'b1000100110101000;
    n11032[81] = 16'b1010001000101010;
    n11032[80] = 16'b0110011011011100;
    n11032[79] = 16'b1110111010110001;
    n11032[78] = 16'b0111011010100100;
    n11032[77] = 16'b0100011001111101;
    n11032[76] = 16'b0001011010000111;
    n11032[75] = 16'b1111101110001011;
    n11032[74] = 16'b1110010111101011;
    n11032[73] = 16'b1011110111000000;
    n11032[72] = 16'b1111110010100011;
    n11032[71] = 16'b1000101100100100;
    n11032[70] = 16'b1110111110111101;
    n11032[69] = 16'b1110011001000001;
    n11032[68] = 16'b0011001100010000;
    n11032[67] = 16'b1110100000111010;
    n11032[66] = 16'b1001011111001111;
    n11032[65] = 16'b0111101010111001;
    n11032[64] = 16'b0101100111110100;
    n11032[63] = 16'b1010110001101110;
    n11032[62] = 16'b1011000100001010;
    n11032[61] = 16'b0101110010000001;
    n11032[60] = 16'b0011111111100001;
    n11032[59] = 16'b0101001101100100;
    n11032[58] = 16'b1101100100001111;
    n11032[57] = 16'b1010100000000010;
    n11032[56] = 16'b0110110001010100;
    n11032[55] = 16'b0111001000111011;
    n11032[54] = 16'b1001110001011100;
    n11032[53] = 16'b0001010000011001;
    n11032[52] = 16'b1001011001101111;
    n11032[51] = 16'b1111101000111110;
    n11032[50] = 16'b1001010111101010;
    n11032[49] = 16'b0000110010110101;
    n11032[48] = 16'b1000010100111111;
    n11032[47] = 16'b0111001101110111;
    n11032[46] = 16'b0001110001000111;
    n11032[45] = 16'b1000111101111111;
    n11032[44] = 16'b0010000111010000;
    n11032[43] = 16'b0111000101101010;
    n11032[42] = 16'b0010010110000100;
    n11032[41] = 16'b0111111000001101;
    n11032[40] = 16'b0100100110010101;
    n11032[39] = 16'b1100001000100011;
    n11032[38] = 16'b1001000000100010;
    n11032[37] = 16'b0011000001110110;
    n11032[36] = 16'b0100100001100110;
    n11032[35] = 16'b0101111110001010;
    n11032[34] = 16'b1100000000011101;
    n11032[33] = 16'b0000010110101100;
    n11032[32] = 16'b0110000101011000;
    n11032[31] = 16'b1100010000110011;
    n11032[30] = 16'b0110111110001110;
    n11032[29] = 16'b0011100100110110;
    n11032[28] = 16'b0000001111000111;
    n11032[27] = 16'b1110010001111001;
    n11032[26] = 16'b1000111011110111;
    n11032[25] = 16'b0111010011011010;
    n11032[24] = 16'b1111111001111000;
    n11032[23] = 16'b1101100000000001;
    n11032[22] = 16'b1011111101011110;
    n11032[21] = 16'b1001101011011000;
    n11032[20] = 16'b0110100010110111;
    n11032[19] = 16'b0010001010111011;
    n11032[18] = 16'b1101011110010010;
    n11032[17] = 16'b0110010011000110;
    n11032[16] = 16'b0011110010011000;
    n11032[15] = 16'b1110001000011111;
    n11032[14] = 16'b1101101010010000;
    n11032[13] = 16'b1010010000100111;
    n11032[12] = 16'b1101000110111110;
    n11032[11] = 16'b0000010000001001;
    n11032[10] = 16'b0110010101010011;
    n11032[9] = 16'b0101011100111001;
    n11032[8] = 16'b0001000010100101;
    n11032[7] = 16'b0110011111011111;
    n11032[6] = 16'b0101100011010110;
    n11032[5] = 16'b1111001011100000;
    n11032[4] = 16'b0011001000010101;
    n11032[3] = 16'b0101110111100110;
    n11032[2] = 16'b0010011111111000;
    n11032[1] = 16'b0010001111000101;
    n11032[0] = 16'b1011000011100011;
    end
  assign n11033_data = n11032[n11027_o];
  /* RTL_PUF/vhdl/random_rom.vhd:275:25  */
endmodule

module ros_selection
  (input  [7:0] challenge,
   input  [255:0] enable,
   output \output );
  (* KEEP="TRUE" *) wire [255:0] sortie_ro;
  (* KEEP="TRUE" *) wire n4873_o;
  (* KEEP="TRUE" *) wire inverseur_n1_ringoscillator_n4874;
  (* KEEP="TRUE" *) wire inverseur_n1_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4877_o;
  (* KEEP="TRUE" *) wire inverseur_n2_ringoscillator_n4878;
  (* KEEP="TRUE" *) wire inverseur_n2_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4881_o;
  (* KEEP="TRUE" *) wire inverseur_n3_ringoscillator_n4882;
  (* KEEP="TRUE" *) wire inverseur_n3_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4885_o;
  (* KEEP="TRUE" *) wire inverseur_n4_ringoscillator_n4886;
  (* KEEP="TRUE" *) wire inverseur_n4_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4889_o;
  (* KEEP="TRUE" *) wire inverseur_n5_ringoscillator_n4890;
  (* KEEP="TRUE" *) wire inverseur_n5_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4893_o;
  (* KEEP="TRUE" *) wire inverseur_n6_ringoscillator_n4894;
  (* KEEP="TRUE" *) wire inverseur_n6_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4897_o;
  (* KEEP="TRUE" *) wire inverseur_n7_ringoscillator_n4898;
  (* KEEP="TRUE" *) wire inverseur_n7_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4901_o;
  (* KEEP="TRUE" *) wire inverseur_n8_ringoscillator_n4902;
  (* KEEP="TRUE" *) wire inverseur_n8_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4905_o;
  (* KEEP="TRUE" *) wire inverseur_n9_ringoscillator_n4906;
  (* KEEP="TRUE" *) wire inverseur_n9_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4909_o;
  (* KEEP="TRUE" *) wire inverseur_n10_ringoscillator_n4910;
  (* KEEP="TRUE" *) wire inverseur_n10_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4913_o;
  (* KEEP="TRUE" *) wire inverseur_n11_ringoscillator_n4914;
  (* KEEP="TRUE" *) wire inverseur_n11_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4917_o;
  (* KEEP="TRUE" *) wire inverseur_n12_ringoscillator_n4918;
  (* KEEP="TRUE" *) wire inverseur_n12_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4921_o;
  (* KEEP="TRUE" *) wire inverseur_n13_ringoscillator_n4922;
  (* KEEP="TRUE" *) wire inverseur_n13_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4925_o;
  (* KEEP="TRUE" *) wire inverseur_n14_ringoscillator_n4926;
  (* KEEP="TRUE" *) wire inverseur_n14_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4929_o;
  (* KEEP="TRUE" *) wire inverseur_n15_ringoscillator_n4930;
  (* KEEP="TRUE" *) wire inverseur_n15_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4933_o;
  (* KEEP="TRUE" *) wire inverseur_n16_ringoscillator_n4934;
  (* KEEP="TRUE" *) wire inverseur_n16_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4937_o;
  (* KEEP="TRUE" *) wire inverseur_n17_ringoscillator_n4938;
  (* KEEP="TRUE" *) wire inverseur_n17_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4941_o;
  (* KEEP="TRUE" *) wire inverseur_n18_ringoscillator_n4942;
  (* KEEP="TRUE" *) wire inverseur_n18_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4945_o;
  (* KEEP="TRUE" *) wire inverseur_n19_ringoscillator_n4946;
  (* KEEP="TRUE" *) wire inverseur_n19_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4949_o;
  (* KEEP="TRUE" *) wire inverseur_n20_ringoscillator_n4950;
  (* KEEP="TRUE" *) wire inverseur_n20_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4953_o;
  (* KEEP="TRUE" *) wire inverseur_n21_ringoscillator_n4954;
  (* KEEP="TRUE" *) wire inverseur_n21_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4957_o;
  (* KEEP="TRUE" *) wire inverseur_n22_ringoscillator_n4958;
  (* KEEP="TRUE" *) wire inverseur_n22_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4961_o;
  (* KEEP="TRUE" *) wire inverseur_n23_ringoscillator_n4962;
  (* KEEP="TRUE" *) wire inverseur_n23_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4965_o;
  (* KEEP="TRUE" *) wire inverseur_n24_ringoscillator_n4966;
  (* KEEP="TRUE" *) wire inverseur_n24_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4969_o;
  (* KEEP="TRUE" *) wire inverseur_n25_ringoscillator_n4970;
  (* KEEP="TRUE" *) wire inverseur_n25_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4973_o;
  (* KEEP="TRUE" *) wire inverseur_n26_ringoscillator_n4974;
  (* KEEP="TRUE" *) wire inverseur_n26_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4977_o;
  (* KEEP="TRUE" *) wire inverseur_n27_ringoscillator_n4978;
  (* KEEP="TRUE" *) wire inverseur_n27_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4981_o;
  (* KEEP="TRUE" *) wire inverseur_n28_ringoscillator_n4982;
  (* KEEP="TRUE" *) wire inverseur_n28_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4985_o;
  (* KEEP="TRUE" *) wire inverseur_n29_ringoscillator_n4986;
  (* KEEP="TRUE" *) wire inverseur_n29_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4989_o;
  (* KEEP="TRUE" *) wire inverseur_n30_ringoscillator_n4990;
  (* KEEP="TRUE" *) wire inverseur_n30_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4993_o;
  (* KEEP="TRUE" *) wire inverseur_n31_ringoscillator_n4994;
  (* KEEP="TRUE" *) wire inverseur_n31_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n4997_o;
  (* KEEP="TRUE" *) wire inverseur_n32_ringoscillator_n4998;
  (* KEEP="TRUE" *) wire inverseur_n32_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5001_o;
  (* KEEP="TRUE" *) wire inverseur_n33_ringoscillator_n5002;
  (* KEEP="TRUE" *) wire inverseur_n33_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5005_o;
  (* KEEP="TRUE" *) wire inverseur_n34_ringoscillator_n5006;
  (* KEEP="TRUE" *) wire inverseur_n34_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5009_o;
  (* KEEP="TRUE" *) wire inverseur_n35_ringoscillator_n5010;
  (* KEEP="TRUE" *) wire inverseur_n35_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5013_o;
  (* KEEP="TRUE" *) wire inverseur_n36_ringoscillator_n5014;
  (* KEEP="TRUE" *) wire inverseur_n36_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5017_o;
  (* KEEP="TRUE" *) wire inverseur_n37_ringoscillator_n5018;
  (* KEEP="TRUE" *) wire inverseur_n37_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5021_o;
  (* KEEP="TRUE" *) wire inverseur_n38_ringoscillator_n5022;
  (* KEEP="TRUE" *) wire inverseur_n38_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5025_o;
  (* KEEP="TRUE" *) wire inverseur_n39_ringoscillator_n5026;
  (* KEEP="TRUE" *) wire inverseur_n39_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5029_o;
  (* KEEP="TRUE" *) wire inverseur_n40_ringoscillator_n5030;
  (* KEEP="TRUE" *) wire inverseur_n40_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5033_o;
  (* KEEP="TRUE" *) wire inverseur_n41_ringoscillator_n5034;
  (* KEEP="TRUE" *) wire inverseur_n41_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5037_o;
  (* KEEP="TRUE" *) wire inverseur_n42_ringoscillator_n5038;
  (* KEEP="TRUE" *) wire inverseur_n42_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5041_o;
  (* KEEP="TRUE" *) wire inverseur_n43_ringoscillator_n5042;
  (* KEEP="TRUE" *) wire inverseur_n43_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5045_o;
  (* KEEP="TRUE" *) wire inverseur_n44_ringoscillator_n5046;
  (* KEEP="TRUE" *) wire inverseur_n44_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5049_o;
  (* KEEP="TRUE" *) wire inverseur_n45_ringoscillator_n5050;
  (* KEEP="TRUE" *) wire inverseur_n45_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5053_o;
  (* KEEP="TRUE" *) wire inverseur_n46_ringoscillator_n5054;
  (* KEEP="TRUE" *) wire inverseur_n46_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5057_o;
  (* KEEP="TRUE" *) wire inverseur_n47_ringoscillator_n5058;
  (* KEEP="TRUE" *) wire inverseur_n47_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5061_o;
  (* KEEP="TRUE" *) wire inverseur_n48_ringoscillator_n5062;
  (* KEEP="TRUE" *) wire inverseur_n48_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5065_o;
  (* KEEP="TRUE" *) wire inverseur_n49_ringoscillator_n5066;
  (* KEEP="TRUE" *) wire inverseur_n49_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5069_o;
  (* KEEP="TRUE" *) wire inverseur_n50_ringoscillator_n5070;
  (* KEEP="TRUE" *) wire inverseur_n50_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5073_o;
  (* KEEP="TRUE" *) wire inverseur_n51_ringoscillator_n5074;
  (* KEEP="TRUE" *) wire inverseur_n51_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5077_o;
  (* KEEP="TRUE" *) wire inverseur_n52_ringoscillator_n5078;
  (* KEEP="TRUE" *) wire inverseur_n52_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5081_o;
  (* KEEP="TRUE" *) wire inverseur_n53_ringoscillator_n5082;
  (* KEEP="TRUE" *) wire inverseur_n53_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5085_o;
  (* KEEP="TRUE" *) wire inverseur_n54_ringoscillator_n5086;
  (* KEEP="TRUE" *) wire inverseur_n54_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5089_o;
  (* KEEP="TRUE" *) wire inverseur_n55_ringoscillator_n5090;
  (* KEEP="TRUE" *) wire inverseur_n55_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5093_o;
  (* KEEP="TRUE" *) wire inverseur_n56_ringoscillator_n5094;
  (* KEEP="TRUE" *) wire inverseur_n56_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5097_o;
  (* KEEP="TRUE" *) wire inverseur_n57_ringoscillator_n5098;
  (* KEEP="TRUE" *) wire inverseur_n57_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5101_o;
  (* KEEP="TRUE" *) wire inverseur_n58_ringoscillator_n5102;
  (* KEEP="TRUE" *) wire inverseur_n58_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5105_o;
  (* KEEP="TRUE" *) wire inverseur_n59_ringoscillator_n5106;
  (* KEEP="TRUE" *) wire inverseur_n59_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5109_o;
  (* KEEP="TRUE" *) wire inverseur_n60_ringoscillator_n5110;
  (* KEEP="TRUE" *) wire inverseur_n60_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5113_o;
  (* KEEP="TRUE" *) wire inverseur_n61_ringoscillator_n5114;
  (* KEEP="TRUE" *) wire inverseur_n61_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5117_o;
  (* KEEP="TRUE" *) wire inverseur_n62_ringoscillator_n5118;
  (* KEEP="TRUE" *) wire inverseur_n62_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5121_o;
  (* KEEP="TRUE" *) wire inverseur_n63_ringoscillator_n5122;
  (* KEEP="TRUE" *) wire inverseur_n63_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5125_o;
  (* KEEP="TRUE" *) wire inverseur_n64_ringoscillator_n5126;
  (* KEEP="TRUE" *) wire inverseur_n64_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5129_o;
  (* KEEP="TRUE" *) wire inverseur_n65_ringoscillator_n5130;
  (* KEEP="TRUE" *) wire inverseur_n65_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5133_o;
  (* KEEP="TRUE" *) wire inverseur_n66_ringoscillator_n5134;
  (* KEEP="TRUE" *) wire inverseur_n66_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5137_o;
  (* KEEP="TRUE" *) wire inverseur_n67_ringoscillator_n5138;
  (* KEEP="TRUE" *) wire inverseur_n67_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5141_o;
  (* KEEP="TRUE" *) wire inverseur_n68_ringoscillator_n5142;
  (* KEEP="TRUE" *) wire inverseur_n68_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5145_o;
  (* KEEP="TRUE" *) wire inverseur_n69_ringoscillator_n5146;
  (* KEEP="TRUE" *) wire inverseur_n69_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5149_o;
  (* KEEP="TRUE" *) wire inverseur_n70_ringoscillator_n5150;
  (* KEEP="TRUE" *) wire inverseur_n70_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5153_o;
  (* KEEP="TRUE" *) wire inverseur_n71_ringoscillator_n5154;
  (* KEEP="TRUE" *) wire inverseur_n71_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5157_o;
  (* KEEP="TRUE" *) wire inverseur_n72_ringoscillator_n5158;
  (* KEEP="TRUE" *) wire inverseur_n72_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5161_o;
  (* KEEP="TRUE" *) wire inverseur_n73_ringoscillator_n5162;
  (* KEEP="TRUE" *) wire inverseur_n73_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5165_o;
  (* KEEP="TRUE" *) wire inverseur_n74_ringoscillator_n5166;
  (* KEEP="TRUE" *) wire inverseur_n74_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5169_o;
  (* KEEP="TRUE" *) wire inverseur_n75_ringoscillator_n5170;
  (* KEEP="TRUE" *) wire inverseur_n75_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5173_o;
  (* KEEP="TRUE" *) wire inverseur_n76_ringoscillator_n5174;
  (* KEEP="TRUE" *) wire inverseur_n76_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5177_o;
  (* KEEP="TRUE" *) wire inverseur_n77_ringoscillator_n5178;
  (* KEEP="TRUE" *) wire inverseur_n77_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5181_o;
  (* KEEP="TRUE" *) wire inverseur_n78_ringoscillator_n5182;
  (* KEEP="TRUE" *) wire inverseur_n78_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5185_o;
  (* KEEP="TRUE" *) wire inverseur_n79_ringoscillator_n5186;
  (* KEEP="TRUE" *) wire inverseur_n79_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5189_o;
  (* KEEP="TRUE" *) wire inverseur_n80_ringoscillator_n5190;
  (* KEEP="TRUE" *) wire inverseur_n80_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5193_o;
  (* KEEP="TRUE" *) wire inverseur_n81_ringoscillator_n5194;
  (* KEEP="TRUE" *) wire inverseur_n81_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5197_o;
  (* KEEP="TRUE" *) wire inverseur_n82_ringoscillator_n5198;
  (* KEEP="TRUE" *) wire inverseur_n82_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5201_o;
  (* KEEP="TRUE" *) wire inverseur_n83_ringoscillator_n5202;
  (* KEEP="TRUE" *) wire inverseur_n83_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5205_o;
  (* KEEP="TRUE" *) wire inverseur_n84_ringoscillator_n5206;
  (* KEEP="TRUE" *) wire inverseur_n84_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5209_o;
  (* KEEP="TRUE" *) wire inverseur_n85_ringoscillator_n5210;
  (* KEEP="TRUE" *) wire inverseur_n85_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5213_o;
  (* KEEP="TRUE" *) wire inverseur_n86_ringoscillator_n5214;
  (* KEEP="TRUE" *) wire inverseur_n86_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5217_o;
  (* KEEP="TRUE" *) wire inverseur_n87_ringoscillator_n5218;
  (* KEEP="TRUE" *) wire inverseur_n87_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5221_o;
  (* KEEP="TRUE" *) wire inverseur_n88_ringoscillator_n5222;
  (* KEEP="TRUE" *) wire inverseur_n88_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5225_o;
  (* KEEP="TRUE" *) wire inverseur_n89_ringoscillator_n5226;
  (* KEEP="TRUE" *) wire inverseur_n89_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5229_o;
  (* KEEP="TRUE" *) wire inverseur_n90_ringoscillator_n5230;
  (* KEEP="TRUE" *) wire inverseur_n90_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5233_o;
  (* KEEP="TRUE" *) wire inverseur_n91_ringoscillator_n5234;
  (* KEEP="TRUE" *) wire inverseur_n91_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5237_o;
  (* KEEP="TRUE" *) wire inverseur_n92_ringoscillator_n5238;
  (* KEEP="TRUE" *) wire inverseur_n92_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5241_o;
  (* KEEP="TRUE" *) wire inverseur_n93_ringoscillator_n5242;
  (* KEEP="TRUE" *) wire inverseur_n93_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5245_o;
  (* KEEP="TRUE" *) wire inverseur_n94_ringoscillator_n5246;
  (* KEEP="TRUE" *) wire inverseur_n94_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5249_o;
  (* KEEP="TRUE" *) wire inverseur_n95_ringoscillator_n5250;
  (* KEEP="TRUE" *) wire inverseur_n95_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5253_o;
  (* KEEP="TRUE" *) wire inverseur_n96_ringoscillator_n5254;
  (* KEEP="TRUE" *) wire inverseur_n96_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5257_o;
  (* KEEP="TRUE" *) wire inverseur_n97_ringoscillator_n5258;
  (* KEEP="TRUE" *) wire inverseur_n97_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5261_o;
  (* KEEP="TRUE" *) wire inverseur_n98_ringoscillator_n5262;
  (* KEEP="TRUE" *) wire inverseur_n98_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5265_o;
  (* KEEP="TRUE" *) wire inverseur_n99_ringoscillator_n5266;
  (* KEEP="TRUE" *) wire inverseur_n99_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5269_o;
  (* KEEP="TRUE" *) wire inverseur_n100_ringoscillator_n5270;
  (* KEEP="TRUE" *) wire inverseur_n100_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5273_o;
  (* KEEP="TRUE" *) wire inverseur_n101_ringoscillator_n5274;
  (* KEEP="TRUE" *) wire inverseur_n101_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5277_o;
  (* KEEP="TRUE" *) wire inverseur_n102_ringoscillator_n5278;
  (* KEEP="TRUE" *) wire inverseur_n102_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5281_o;
  (* KEEP="TRUE" *) wire inverseur_n103_ringoscillator_n5282;
  (* KEEP="TRUE" *) wire inverseur_n103_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5285_o;
  (* KEEP="TRUE" *) wire inverseur_n104_ringoscillator_n5286;
  (* KEEP="TRUE" *) wire inverseur_n104_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5289_o;
  (* KEEP="TRUE" *) wire inverseur_n105_ringoscillator_n5290;
  (* KEEP="TRUE" *) wire inverseur_n105_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5293_o;
  (* KEEP="TRUE" *) wire inverseur_n106_ringoscillator_n5294;
  (* KEEP="TRUE" *) wire inverseur_n106_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5297_o;
  (* KEEP="TRUE" *) wire inverseur_n107_ringoscillator_n5298;
  (* KEEP="TRUE" *) wire inverseur_n107_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5301_o;
  (* KEEP="TRUE" *) wire inverseur_n108_ringoscillator_n5302;
  (* KEEP="TRUE" *) wire inverseur_n108_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5305_o;
  (* KEEP="TRUE" *) wire inverseur_n109_ringoscillator_n5306;
  (* KEEP="TRUE" *) wire inverseur_n109_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5309_o;
  (* KEEP="TRUE" *) wire inverseur_n110_ringoscillator_n5310;
  (* KEEP="TRUE" *) wire inverseur_n110_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5313_o;
  (* KEEP="TRUE" *) wire inverseur_n111_ringoscillator_n5314;
  (* KEEP="TRUE" *) wire inverseur_n111_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5317_o;
  (* KEEP="TRUE" *) wire inverseur_n112_ringoscillator_n5318;
  (* KEEP="TRUE" *) wire inverseur_n112_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5321_o;
  (* KEEP="TRUE" *) wire inverseur_n113_ringoscillator_n5322;
  (* KEEP="TRUE" *) wire inverseur_n113_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5325_o;
  (* KEEP="TRUE" *) wire inverseur_n114_ringoscillator_n5326;
  (* KEEP="TRUE" *) wire inverseur_n114_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5329_o;
  (* KEEP="TRUE" *) wire inverseur_n115_ringoscillator_n5330;
  (* KEEP="TRUE" *) wire inverseur_n115_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5333_o;
  (* KEEP="TRUE" *) wire inverseur_n116_ringoscillator_n5334;
  (* KEEP="TRUE" *) wire inverseur_n116_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5337_o;
  (* KEEP="TRUE" *) wire inverseur_n117_ringoscillator_n5338;
  (* KEEP="TRUE" *) wire inverseur_n117_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5341_o;
  (* KEEP="TRUE" *) wire inverseur_n118_ringoscillator_n5342;
  (* KEEP="TRUE" *) wire inverseur_n118_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5345_o;
  (* KEEP="TRUE" *) wire inverseur_n119_ringoscillator_n5346;
  (* KEEP="TRUE" *) wire inverseur_n119_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5349_o;
  (* KEEP="TRUE" *) wire inverseur_n120_ringoscillator_n5350;
  (* KEEP="TRUE" *) wire inverseur_n120_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5353_o;
  (* KEEP="TRUE" *) wire inverseur_n121_ringoscillator_n5354;
  (* KEEP="TRUE" *) wire inverseur_n121_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5357_o;
  (* KEEP="TRUE" *) wire inverseur_n122_ringoscillator_n5358;
  (* KEEP="TRUE" *) wire inverseur_n122_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5361_o;
  (* KEEP="TRUE" *) wire inverseur_n123_ringoscillator_n5362;
  (* KEEP="TRUE" *) wire inverseur_n123_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5365_o;
  (* KEEP="TRUE" *) wire inverseur_n124_ringoscillator_n5366;
  (* KEEP="TRUE" *) wire inverseur_n124_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5369_o;
  (* KEEP="TRUE" *) wire inverseur_n125_ringoscillator_n5370;
  (* KEEP="TRUE" *) wire inverseur_n125_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5373_o;
  (* KEEP="TRUE" *) wire inverseur_n126_ringoscillator_n5374;
  (* KEEP="TRUE" *) wire inverseur_n126_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5377_o;
  (* KEEP="TRUE" *) wire inverseur_n127_ringoscillator_n5378;
  (* KEEP="TRUE" *) wire inverseur_n127_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5381_o;
  (* KEEP="TRUE" *) wire inverseur_n128_ringoscillator_n5382;
  (* KEEP="TRUE" *) wire inverseur_n128_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5385_o;
  (* KEEP="TRUE" *) wire inverseur_n129_ringoscillator_n5386;
  (* KEEP="TRUE" *) wire inverseur_n129_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5389_o;
  (* KEEP="TRUE" *) wire inverseur_n130_ringoscillator_n5390;
  (* KEEP="TRUE" *) wire inverseur_n130_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5393_o;
  (* KEEP="TRUE" *) wire inverseur_n131_ringoscillator_n5394;
  (* KEEP="TRUE" *) wire inverseur_n131_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5397_o;
  (* KEEP="TRUE" *) wire inverseur_n132_ringoscillator_n5398;
  (* KEEP="TRUE" *) wire inverseur_n132_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5401_o;
  (* KEEP="TRUE" *) wire inverseur_n133_ringoscillator_n5402;
  (* KEEP="TRUE" *) wire inverseur_n133_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5405_o;
  (* KEEP="TRUE" *) wire inverseur_n134_ringoscillator_n5406;
  (* KEEP="TRUE" *) wire inverseur_n134_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5409_o;
  (* KEEP="TRUE" *) wire inverseur_n135_ringoscillator_n5410;
  (* KEEP="TRUE" *) wire inverseur_n135_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5413_o;
  (* KEEP="TRUE" *) wire inverseur_n136_ringoscillator_n5414;
  (* KEEP="TRUE" *) wire inverseur_n136_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5417_o;
  (* KEEP="TRUE" *) wire inverseur_n137_ringoscillator_n5418;
  (* KEEP="TRUE" *) wire inverseur_n137_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5421_o;
  (* KEEP="TRUE" *) wire inverseur_n138_ringoscillator_n5422;
  (* KEEP="TRUE" *) wire inverseur_n138_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5425_o;
  (* KEEP="TRUE" *) wire inverseur_n139_ringoscillator_n5426;
  (* KEEP="TRUE" *) wire inverseur_n139_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5429_o;
  (* KEEP="TRUE" *) wire inverseur_n140_ringoscillator_n5430;
  (* KEEP="TRUE" *) wire inverseur_n140_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5433_o;
  (* KEEP="TRUE" *) wire inverseur_n141_ringoscillator_n5434;
  (* KEEP="TRUE" *) wire inverseur_n141_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5437_o;
  (* KEEP="TRUE" *) wire inverseur_n142_ringoscillator_n5438;
  (* KEEP="TRUE" *) wire inverseur_n142_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5441_o;
  (* KEEP="TRUE" *) wire inverseur_n143_ringoscillator_n5442;
  (* KEEP="TRUE" *) wire inverseur_n143_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5445_o;
  (* KEEP="TRUE" *) wire inverseur_n144_ringoscillator_n5446;
  (* KEEP="TRUE" *) wire inverseur_n144_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5449_o;
  (* KEEP="TRUE" *) wire inverseur_n145_ringoscillator_n5450;
  (* KEEP="TRUE" *) wire inverseur_n145_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5453_o;
  (* KEEP="TRUE" *) wire inverseur_n146_ringoscillator_n5454;
  (* KEEP="TRUE" *) wire inverseur_n146_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5457_o;
  (* KEEP="TRUE" *) wire inverseur_n147_ringoscillator_n5458;
  (* KEEP="TRUE" *) wire inverseur_n147_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5461_o;
  (* KEEP="TRUE" *) wire inverseur_n148_ringoscillator_n5462;
  (* KEEP="TRUE" *) wire inverseur_n148_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5465_o;
  (* KEEP="TRUE" *) wire inverseur_n149_ringoscillator_n5466;
  (* KEEP="TRUE" *) wire inverseur_n149_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5469_o;
  (* KEEP="TRUE" *) wire inverseur_n150_ringoscillator_n5470;
  (* KEEP="TRUE" *) wire inverseur_n150_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5473_o;
  (* KEEP="TRUE" *) wire inverseur_n151_ringoscillator_n5474;
  (* KEEP="TRUE" *) wire inverseur_n151_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5477_o;
  (* KEEP="TRUE" *) wire inverseur_n152_ringoscillator_n5478;
  (* KEEP="TRUE" *) wire inverseur_n152_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5481_o;
  (* KEEP="TRUE" *) wire inverseur_n153_ringoscillator_n5482;
  (* KEEP="TRUE" *) wire inverseur_n153_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5485_o;
  (* KEEP="TRUE" *) wire inverseur_n154_ringoscillator_n5486;
  (* KEEP="TRUE" *) wire inverseur_n154_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5489_o;
  (* KEEP="TRUE" *) wire inverseur_n155_ringoscillator_n5490;
  (* KEEP="TRUE" *) wire inverseur_n155_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5493_o;
  (* KEEP="TRUE" *) wire inverseur_n156_ringoscillator_n5494;
  (* KEEP="TRUE" *) wire inverseur_n156_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5497_o;
  (* KEEP="TRUE" *) wire inverseur_n157_ringoscillator_n5498;
  (* KEEP="TRUE" *) wire inverseur_n157_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5501_o;
  (* KEEP="TRUE" *) wire inverseur_n158_ringoscillator_n5502;
  (* KEEP="TRUE" *) wire inverseur_n158_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5505_o;
  (* KEEP="TRUE" *) wire inverseur_n159_ringoscillator_n5506;
  (* KEEP="TRUE" *) wire inverseur_n159_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5509_o;
  (* KEEP="TRUE" *) wire inverseur_n160_ringoscillator_n5510;
  (* KEEP="TRUE" *) wire inverseur_n160_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5513_o;
  (* KEEP="TRUE" *) wire inverseur_n161_ringoscillator_n5514;
  (* KEEP="TRUE" *) wire inverseur_n161_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5517_o;
  (* KEEP="TRUE" *) wire inverseur_n162_ringoscillator_n5518;
  (* KEEP="TRUE" *) wire inverseur_n162_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5521_o;
  (* KEEP="TRUE" *) wire inverseur_n163_ringoscillator_n5522;
  (* KEEP="TRUE" *) wire inverseur_n163_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5525_o;
  (* KEEP="TRUE" *) wire inverseur_n164_ringoscillator_n5526;
  (* KEEP="TRUE" *) wire inverseur_n164_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5529_o;
  (* KEEP="TRUE" *) wire inverseur_n165_ringoscillator_n5530;
  (* KEEP="TRUE" *) wire inverseur_n165_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5533_o;
  (* KEEP="TRUE" *) wire inverseur_n166_ringoscillator_n5534;
  (* KEEP="TRUE" *) wire inverseur_n166_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5537_o;
  (* KEEP="TRUE" *) wire inverseur_n167_ringoscillator_n5538;
  (* KEEP="TRUE" *) wire inverseur_n167_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5541_o;
  (* KEEP="TRUE" *) wire inverseur_n168_ringoscillator_n5542;
  (* KEEP="TRUE" *) wire inverseur_n168_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5545_o;
  (* KEEP="TRUE" *) wire inverseur_n169_ringoscillator_n5546;
  (* KEEP="TRUE" *) wire inverseur_n169_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5549_o;
  (* KEEP="TRUE" *) wire inverseur_n170_ringoscillator_n5550;
  (* KEEP="TRUE" *) wire inverseur_n170_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5553_o;
  (* KEEP="TRUE" *) wire inverseur_n171_ringoscillator_n5554;
  (* KEEP="TRUE" *) wire inverseur_n171_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5557_o;
  (* KEEP="TRUE" *) wire inverseur_n172_ringoscillator_n5558;
  (* KEEP="TRUE" *) wire inverseur_n172_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5561_o;
  (* KEEP="TRUE" *) wire inverseur_n173_ringoscillator_n5562;
  (* KEEP="TRUE" *) wire inverseur_n173_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5565_o;
  (* KEEP="TRUE" *) wire inverseur_n174_ringoscillator_n5566;
  (* KEEP="TRUE" *) wire inverseur_n174_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5569_o;
  (* KEEP="TRUE" *) wire inverseur_n175_ringoscillator_n5570;
  (* KEEP="TRUE" *) wire inverseur_n175_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5573_o;
  (* KEEP="TRUE" *) wire inverseur_n176_ringoscillator_n5574;
  (* KEEP="TRUE" *) wire inverseur_n176_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5577_o;
  (* KEEP="TRUE" *) wire inverseur_n177_ringoscillator_n5578;
  (* KEEP="TRUE" *) wire inverseur_n177_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5581_o;
  (* KEEP="TRUE" *) wire inverseur_n178_ringoscillator_n5582;
  (* KEEP="TRUE" *) wire inverseur_n178_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5585_o;
  (* KEEP="TRUE" *) wire inverseur_n179_ringoscillator_n5586;
  (* KEEP="TRUE" *) wire inverseur_n179_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5589_o;
  (* KEEP="TRUE" *) wire inverseur_n180_ringoscillator_n5590;
  (* KEEP="TRUE" *) wire inverseur_n180_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5593_o;
  (* KEEP="TRUE" *) wire inverseur_n181_ringoscillator_n5594;
  (* KEEP="TRUE" *) wire inverseur_n181_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5597_o;
  (* KEEP="TRUE" *) wire inverseur_n182_ringoscillator_n5598;
  (* KEEP="TRUE" *) wire inverseur_n182_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5601_o;
  (* KEEP="TRUE" *) wire inverseur_n183_ringoscillator_n5602;
  (* KEEP="TRUE" *) wire inverseur_n183_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5605_o;
  (* KEEP="TRUE" *) wire inverseur_n184_ringoscillator_n5606;
  (* KEEP="TRUE" *) wire inverseur_n184_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5609_o;
  (* KEEP="TRUE" *) wire inverseur_n185_ringoscillator_n5610;
  (* KEEP="TRUE" *) wire inverseur_n185_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5613_o;
  (* KEEP="TRUE" *) wire inverseur_n186_ringoscillator_n5614;
  (* KEEP="TRUE" *) wire inverseur_n186_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5617_o;
  (* KEEP="TRUE" *) wire inverseur_n187_ringoscillator_n5618;
  (* KEEP="TRUE" *) wire inverseur_n187_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5621_o;
  (* KEEP="TRUE" *) wire inverseur_n188_ringoscillator_n5622;
  (* KEEP="TRUE" *) wire inverseur_n188_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5625_o;
  (* KEEP="TRUE" *) wire inverseur_n189_ringoscillator_n5626;
  (* KEEP="TRUE" *) wire inverseur_n189_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5629_o;
  (* KEEP="TRUE" *) wire inverseur_n190_ringoscillator_n5630;
  (* KEEP="TRUE" *) wire inverseur_n190_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5633_o;
  (* KEEP="TRUE" *) wire inverseur_n191_ringoscillator_n5634;
  (* KEEP="TRUE" *) wire inverseur_n191_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5637_o;
  (* KEEP="TRUE" *) wire inverseur_n192_ringoscillator_n5638;
  (* KEEP="TRUE" *) wire inverseur_n192_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5641_o;
  (* KEEP="TRUE" *) wire inverseur_n193_ringoscillator_n5642;
  (* KEEP="TRUE" *) wire inverseur_n193_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5645_o;
  (* KEEP="TRUE" *) wire inverseur_n194_ringoscillator_n5646;
  (* KEEP="TRUE" *) wire inverseur_n194_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5649_o;
  (* KEEP="TRUE" *) wire inverseur_n195_ringoscillator_n5650;
  (* KEEP="TRUE" *) wire inverseur_n195_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5653_o;
  (* KEEP="TRUE" *) wire inverseur_n196_ringoscillator_n5654;
  (* KEEP="TRUE" *) wire inverseur_n196_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5657_o;
  (* KEEP="TRUE" *) wire inverseur_n197_ringoscillator_n5658;
  (* KEEP="TRUE" *) wire inverseur_n197_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5661_o;
  (* KEEP="TRUE" *) wire inverseur_n198_ringoscillator_n5662;
  (* KEEP="TRUE" *) wire inverseur_n198_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5665_o;
  (* KEEP="TRUE" *) wire inverseur_n199_ringoscillator_n5666;
  (* KEEP="TRUE" *) wire inverseur_n199_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5669_o;
  (* KEEP="TRUE" *) wire inverseur_n200_ringoscillator_n5670;
  (* KEEP="TRUE" *) wire inverseur_n200_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5673_o;
  (* KEEP="TRUE" *) wire inverseur_n201_ringoscillator_n5674;
  (* KEEP="TRUE" *) wire inverseur_n201_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5677_o;
  (* KEEP="TRUE" *) wire inverseur_n202_ringoscillator_n5678;
  (* KEEP="TRUE" *) wire inverseur_n202_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5681_o;
  (* KEEP="TRUE" *) wire inverseur_n203_ringoscillator_n5682;
  (* KEEP="TRUE" *) wire inverseur_n203_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5685_o;
  (* KEEP="TRUE" *) wire inverseur_n204_ringoscillator_n5686;
  (* KEEP="TRUE" *) wire inverseur_n204_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5689_o;
  (* KEEP="TRUE" *) wire inverseur_n205_ringoscillator_n5690;
  (* KEEP="TRUE" *) wire inverseur_n205_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5693_o;
  (* KEEP="TRUE" *) wire inverseur_n206_ringoscillator_n5694;
  (* KEEP="TRUE" *) wire inverseur_n206_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5697_o;
  (* KEEP="TRUE" *) wire inverseur_n207_ringoscillator_n5698;
  (* KEEP="TRUE" *) wire inverseur_n207_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5701_o;
  (* KEEP="TRUE" *) wire inverseur_n208_ringoscillator_n5702;
  (* KEEP="TRUE" *) wire inverseur_n208_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5705_o;
  (* KEEP="TRUE" *) wire inverseur_n209_ringoscillator_n5706;
  (* KEEP="TRUE" *) wire inverseur_n209_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5709_o;
  (* KEEP="TRUE" *) wire inverseur_n210_ringoscillator_n5710;
  (* KEEP="TRUE" *) wire inverseur_n210_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5713_o;
  (* KEEP="TRUE" *) wire inverseur_n211_ringoscillator_n5714;
  (* KEEP="TRUE" *) wire inverseur_n211_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5717_o;
  (* KEEP="TRUE" *) wire inverseur_n212_ringoscillator_n5718;
  (* KEEP="TRUE" *) wire inverseur_n212_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5721_o;
  (* KEEP="TRUE" *) wire inverseur_n213_ringoscillator_n5722;
  (* KEEP="TRUE" *) wire inverseur_n213_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5725_o;
  (* KEEP="TRUE" *) wire inverseur_n214_ringoscillator_n5726;
  (* KEEP="TRUE" *) wire inverseur_n214_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5729_o;
  (* KEEP="TRUE" *) wire inverseur_n215_ringoscillator_n5730;
  (* KEEP="TRUE" *) wire inverseur_n215_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5733_o;
  (* KEEP="TRUE" *) wire inverseur_n216_ringoscillator_n5734;
  (* KEEP="TRUE" *) wire inverseur_n216_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5737_o;
  (* KEEP="TRUE" *) wire inverseur_n217_ringoscillator_n5738;
  (* KEEP="TRUE" *) wire inverseur_n217_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5741_o;
  (* KEEP="TRUE" *) wire inverseur_n218_ringoscillator_n5742;
  (* KEEP="TRUE" *) wire inverseur_n218_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5745_o;
  (* KEEP="TRUE" *) wire inverseur_n219_ringoscillator_n5746;
  (* KEEP="TRUE" *) wire inverseur_n219_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5749_o;
  (* KEEP="TRUE" *) wire inverseur_n220_ringoscillator_n5750;
  (* KEEP="TRUE" *) wire inverseur_n220_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5753_o;
  (* KEEP="TRUE" *) wire inverseur_n221_ringoscillator_n5754;
  (* KEEP="TRUE" *) wire inverseur_n221_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5757_o;
  (* KEEP="TRUE" *) wire inverseur_n222_ringoscillator_n5758;
  (* KEEP="TRUE" *) wire inverseur_n222_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5761_o;
  (* KEEP="TRUE" *) wire inverseur_n223_ringoscillator_n5762;
  (* KEEP="TRUE" *) wire inverseur_n223_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5765_o;
  (* KEEP="TRUE" *) wire inverseur_n224_ringoscillator_n5766;
  (* KEEP="TRUE" *) wire inverseur_n224_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5769_o;
  (* KEEP="TRUE" *) wire inverseur_n225_ringoscillator_n5770;
  (* KEEP="TRUE" *) wire inverseur_n225_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5773_o;
  (* KEEP="TRUE" *) wire inverseur_n226_ringoscillator_n5774;
  (* KEEP="TRUE" *) wire inverseur_n226_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5777_o;
  (* KEEP="TRUE" *) wire inverseur_n227_ringoscillator_n5778;
  (* KEEP="TRUE" *) wire inverseur_n227_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5781_o;
  (* KEEP="TRUE" *) wire inverseur_n228_ringoscillator_n5782;
  (* KEEP="TRUE" *) wire inverseur_n228_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5785_o;
  (* KEEP="TRUE" *) wire inverseur_n229_ringoscillator_n5786;
  (* KEEP="TRUE" *) wire inverseur_n229_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5789_o;
  (* KEEP="TRUE" *) wire inverseur_n230_ringoscillator_n5790;
  (* KEEP="TRUE" *) wire inverseur_n230_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5793_o;
  (* KEEP="TRUE" *) wire inverseur_n231_ringoscillator_n5794;
  (* KEEP="TRUE" *) wire inverseur_n231_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5797_o;
  (* KEEP="TRUE" *) wire inverseur_n232_ringoscillator_n5798;
  (* KEEP="TRUE" *) wire inverseur_n232_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5801_o;
  (* KEEP="TRUE" *) wire inverseur_n233_ringoscillator_n5802;
  (* KEEP="TRUE" *) wire inverseur_n233_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5805_o;
  (* KEEP="TRUE" *) wire inverseur_n234_ringoscillator_n5806;
  (* KEEP="TRUE" *) wire inverseur_n234_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5809_o;
  (* KEEP="TRUE" *) wire inverseur_n235_ringoscillator_n5810;
  (* KEEP="TRUE" *) wire inverseur_n235_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5813_o;
  (* KEEP="TRUE" *) wire inverseur_n236_ringoscillator_n5814;
  (* KEEP="TRUE" *) wire inverseur_n236_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5817_o;
  (* KEEP="TRUE" *) wire inverseur_n237_ringoscillator_n5818;
  (* KEEP="TRUE" *) wire inverseur_n237_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5821_o;
  (* KEEP="TRUE" *) wire inverseur_n238_ringoscillator_n5822;
  (* KEEP="TRUE" *) wire inverseur_n238_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5825_o;
  (* KEEP="TRUE" *) wire inverseur_n239_ringoscillator_n5826;
  (* KEEP="TRUE" *) wire inverseur_n239_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5829_o;
  (* KEEP="TRUE" *) wire inverseur_n240_ringoscillator_n5830;
  (* KEEP="TRUE" *) wire inverseur_n240_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5833_o;
  (* KEEP="TRUE" *) wire inverseur_n241_ringoscillator_n5834;
  (* KEEP="TRUE" *) wire inverseur_n241_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5837_o;
  (* KEEP="TRUE" *) wire inverseur_n242_ringoscillator_n5838;
  (* KEEP="TRUE" *) wire inverseur_n242_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5841_o;
  (* KEEP="TRUE" *) wire inverseur_n243_ringoscillator_n5842;
  (* KEEP="TRUE" *) wire inverseur_n243_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5845_o;
  (* KEEP="TRUE" *) wire inverseur_n244_ringoscillator_n5846;
  (* KEEP="TRUE" *) wire inverseur_n244_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5849_o;
  (* KEEP="TRUE" *) wire inverseur_n245_ringoscillator_n5850;
  (* KEEP="TRUE" *) wire inverseur_n245_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5853_o;
  (* KEEP="TRUE" *) wire inverseur_n246_ringoscillator_n5854;
  (* KEEP="TRUE" *) wire inverseur_n246_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5857_o;
  (* KEEP="TRUE" *) wire inverseur_n247_ringoscillator_n5858;
  (* KEEP="TRUE" *) wire inverseur_n247_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5861_o;
  (* KEEP="TRUE" *) wire inverseur_n248_ringoscillator_n5862;
  (* KEEP="TRUE" *) wire inverseur_n248_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5865_o;
  (* KEEP="TRUE" *) wire inverseur_n249_ringoscillator_n5866;
  (* KEEP="TRUE" *) wire inverseur_n249_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5869_o;
  (* KEEP="TRUE" *) wire inverseur_n250_ringoscillator_n5870;
  (* KEEP="TRUE" *) wire inverseur_n250_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5873_o;
  (* KEEP="TRUE" *) wire inverseur_n251_ringoscillator_n5874;
  (* KEEP="TRUE" *) wire inverseur_n251_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5877_o;
  (* KEEP="TRUE" *) wire inverseur_n252_ringoscillator_n5878;
  (* KEEP="TRUE" *) wire inverseur_n252_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5881_o;
  (* KEEP="TRUE" *) wire inverseur_n253_ringoscillator_n5882;
  (* KEEP="TRUE" *) wire inverseur_n253_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5885_o;
  (* KEEP="TRUE" *) wire inverseur_n254_ringoscillator_n5886;
  (* KEEP="TRUE" *) wire inverseur_n254_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5889_o;
  (* KEEP="TRUE" *) wire inverseur_n255_ringoscillator_n5890;
  (* KEEP="TRUE" *) wire inverseur_n255_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5893_o;
  (* KEEP="TRUE" *) wire inverseur_n256_ringoscillator_n5894;
  (* KEEP="TRUE" *) wire inverseur_n256_ringoscillator_ro_out;
  (* KEEP="TRUE" *) wire n5902_o;
  (* KEEP="TRUE" *) wire n5903_o;
  (* KEEP="TRUE" *) wire n5913_o;
  (* KEEP="TRUE" *) wire n5916_o;
  (* KEEP="TRUE" *) wire n5917_o;
  (* KEEP="TRUE" *) wire n5918_o;
  (* KEEP="TRUE" *) wire n5920_o;
  (* KEEP="TRUE" *) wire n5924_o;
  (* KEEP="TRUE" *) wire n5925_o;
  (* KEEP="TRUE" *) wire n5927_o;
  (* KEEP="TRUE" *) wire n5928_o;
  (* KEEP="TRUE" *) wire n5929_o;
  (* KEEP="TRUE" *) wire n5931_o;
  (* KEEP="TRUE" *) wire n5932_o;
  (* KEEP="TRUE" *) wire n5934_o;
  (* KEEP="TRUE" *) wire n5935_o;
  (* KEEP="TRUE" *) wire n5936_o;
  (* KEEP="TRUE" *) wire n5938_o;
  (* KEEP="TRUE" *) wire n5942_o;
  (* KEEP="TRUE" *) wire n5943_o;
  (* KEEP="TRUE" *) wire n5945_o;
  (* KEEP="TRUE" *) wire n5946_o;
  (* KEEP="TRUE" *) wire n5947_o;
  (* KEEP="TRUE" *) wire n5949_o;
  (* KEEP="TRUE" *) wire n5950_o;
  (* KEEP="TRUE" *) wire n5952_o;
  (* KEEP="TRUE" *) wire n5953_o;
  (* KEEP="TRUE" *) wire n5954_o;
  (* KEEP="TRUE" *) wire n5956_o;
  (* KEEP="TRUE" *) wire n5960_o;
  (* KEEP="TRUE" *) wire n5961_o;
  (* KEEP="TRUE" *) wire n5963_o;
  (* KEEP="TRUE" *) wire n5964_o;
  (* KEEP="TRUE" *) wire n5965_o;
  (* KEEP="TRUE" *) wire n5967_o;
  (* KEEP="TRUE" *) wire n5968_o;
  (* KEEP="TRUE" *) wire n5970_o;
  (* KEEP="TRUE" *) wire n5971_o;
  (* KEEP="TRUE" *) wire n5972_o;
  (* KEEP="TRUE" *) wire n5974_o;
  (* KEEP="TRUE" *) wire n5978_o;
  (* KEEP="TRUE" *) wire n5979_o;
  (* KEEP="TRUE" *) wire n5981_o;
  (* KEEP="TRUE" *) wire n5982_o;
  (* KEEP="TRUE" *) wire n5983_o;
  (* KEEP="TRUE" *) wire n5985_o;
  (* KEEP="TRUE" *) wire n5986_o;
  (* KEEP="TRUE" *) wire n5988_o;
  (* KEEP="TRUE" *) wire n5989_o;
  (* KEEP="TRUE" *) wire n5990_o;
  (* KEEP="TRUE" *) wire n5992_o;
  (* KEEP="TRUE" *) wire n5996_o;
  (* KEEP="TRUE" *) wire n5997_o;
  (* KEEP="TRUE" *) wire n5999_o;
  (* KEEP="TRUE" *) wire n6000_o;
  (* KEEP="TRUE" *) wire n6001_o;
  (* KEEP="TRUE" *) wire n6003_o;
  (* KEEP="TRUE" *) wire n6004_o;
  (* KEEP="TRUE" *) wire n6006_o;
  (* KEEP="TRUE" *) wire n6007_o;
  (* KEEP="TRUE" *) wire n6008_o;
  (* KEEP="TRUE" *) wire n6010_o;
  (* KEEP="TRUE" *) wire n6014_o;
  (* KEEP="TRUE" *) wire n6015_o;
  (* KEEP="TRUE" *) wire n6017_o;
  (* KEEP="TRUE" *) wire n6018_o;
  (* KEEP="TRUE" *) wire n6019_o;
  (* KEEP="TRUE" *) wire n6021_o;
  (* KEEP="TRUE" *) wire n6022_o;
  (* KEEP="TRUE" *) wire n6024_o;
  (* KEEP="TRUE" *) wire n6025_o;
  (* KEEP="TRUE" *) wire n6026_o;
  (* KEEP="TRUE" *) wire n6028_o;
  (* KEEP="TRUE" *) wire n6032_o;
  (* KEEP="TRUE" *) wire n6033_o;
  (* KEEP="TRUE" *) wire n6035_o;
  (* KEEP="TRUE" *) wire n6036_o;
  (* KEEP="TRUE" *) wire n6037_o;
  (* KEEP="TRUE" *) wire n6039_o;
  (* KEEP="TRUE" *) wire n6040_o;
  (* KEEP="TRUE" *) wire n6042_o;
  (* KEEP="TRUE" *) wire n6043_o;
  (* KEEP="TRUE" *) wire n6044_o;
  (* KEEP="TRUE" *) wire n6046_o;
  (* KEEP="TRUE" *) wire n6050_o;
  (* KEEP="TRUE" *) wire n6051_o;
  (* KEEP="TRUE" *) wire n6053_o;
  (* KEEP="TRUE" *) wire n6054_o;
  (* KEEP="TRUE" *) wire n6055_o;
  (* KEEP="TRUE" *) wire n6057_o;
  (* KEEP="TRUE" *) wire n6058_o;
  (* KEEP="TRUE" *) wire n6060_o;
  (* KEEP="TRUE" *) wire n6061_o;
  (* KEEP="TRUE" *) wire n6062_o;
  (* KEEP="TRUE" *) wire n6064_o;
  (* KEEP="TRUE" *) wire n6068_o;
  (* KEEP="TRUE" *) wire n6069_o;
  (* KEEP="TRUE" *) wire n6071_o;
  (* KEEP="TRUE" *) wire n6072_o;
  (* KEEP="TRUE" *) wire n6073_o;
  (* KEEP="TRUE" *) wire n6075_o;
  (* KEEP="TRUE" *) wire n6076_o;
  (* KEEP="TRUE" *) wire n6078_o;
  (* KEEP="TRUE" *) wire n6079_o;
  (* KEEP="TRUE" *) wire n6080_o;
  (* KEEP="TRUE" *) wire n6082_o;
  (* KEEP="TRUE" *) wire n6086_o;
  (* KEEP="TRUE" *) wire n6087_o;
  (* KEEP="TRUE" *) wire n6089_o;
  (* KEEP="TRUE" *) wire n6090_o;
  (* KEEP="TRUE" *) wire n6091_o;
  (* KEEP="TRUE" *) wire n6093_o;
  (* KEEP="TRUE" *) wire n6094_o;
  (* KEEP="TRUE" *) wire n6096_o;
  (* KEEP="TRUE" *) wire n6097_o;
  (* KEEP="TRUE" *) wire n6098_o;
  (* KEEP="TRUE" *) wire n6100_o;
  (* KEEP="TRUE" *) wire n6104_o;
  (* KEEP="TRUE" *) wire n6105_o;
  (* KEEP="TRUE" *) wire n6107_o;
  (* KEEP="TRUE" *) wire n6108_o;
  (* KEEP="TRUE" *) wire n6109_o;
  (* KEEP="TRUE" *) wire n6111_o;
  (* KEEP="TRUE" *) wire n6112_o;
  (* KEEP="TRUE" *) wire n6114_o;
  (* KEEP="TRUE" *) wire n6115_o;
  (* KEEP="TRUE" *) wire n6116_o;
  (* KEEP="TRUE" *) wire n6118_o;
  (* KEEP="TRUE" *) wire n6122_o;
  (* KEEP="TRUE" *) wire n6123_o;
  (* KEEP="TRUE" *) wire n6125_o;
  (* KEEP="TRUE" *) wire n6126_o;
  (* KEEP="TRUE" *) wire n6127_o;
  (* KEEP="TRUE" *) wire n6129_o;
  (* KEEP="TRUE" *) wire n6130_o;
  (* KEEP="TRUE" *) wire n6132_o;
  (* KEEP="TRUE" *) wire n6133_o;
  (* KEEP="TRUE" *) wire n6134_o;
  (* KEEP="TRUE" *) wire n6136_o;
  (* KEEP="TRUE" *) wire n6140_o;
  (* KEEP="TRUE" *) wire n6141_o;
  (* KEEP="TRUE" *) wire n6143_o;
  (* KEEP="TRUE" *) wire n6144_o;
  (* KEEP="TRUE" *) wire n6145_o;
  (* KEEP="TRUE" *) wire n6147_o;
  (* KEEP="TRUE" *) wire n6148_o;
  (* KEEP="TRUE" *) wire n6150_o;
  (* KEEP="TRUE" *) wire n6151_o;
  (* KEEP="TRUE" *) wire n6152_o;
  (* KEEP="TRUE" *) wire n6154_o;
  (* KEEP="TRUE" *) wire n6158_o;
  (* KEEP="TRUE" *) wire n6159_o;
  (* KEEP="TRUE" *) wire n6161_o;
  (* KEEP="TRUE" *) wire n6162_o;
  (* KEEP="TRUE" *) wire n6163_o;
  (* KEEP="TRUE" *) wire n6165_o;
  (* KEEP="TRUE" *) wire n6166_o;
  (* KEEP="TRUE" *) wire n6168_o;
  (* KEEP="TRUE" *) wire n6169_o;
  (* KEEP="TRUE" *) wire n6170_o;
  (* KEEP="TRUE" *) wire n6172_o;
  (* KEEP="TRUE" *) wire n6176_o;
  (* KEEP="TRUE" *) wire n6177_o;
  (* KEEP="TRUE" *) wire n6179_o;
  (* KEEP="TRUE" *) wire n6180_o;
  (* KEEP="TRUE" *) wire n6181_o;
  (* KEEP="TRUE" *) wire n6183_o;
  (* KEEP="TRUE" *) wire n6184_o;
  (* KEEP="TRUE" *) wire n6186_o;
  (* KEEP="TRUE" *) wire n6187_o;
  (* KEEP="TRUE" *) wire n6188_o;
  (* KEEP="TRUE" *) wire n6190_o;
  (* KEEP="TRUE" *) wire n6194_o;
  (* KEEP="TRUE" *) wire n6195_o;
  (* KEEP="TRUE" *) wire n6197_o;
  (* KEEP="TRUE" *) wire n6198_o;
  (* KEEP="TRUE" *) wire n6199_o;
  (* KEEP="TRUE" *) wire n6201_o;
  (* KEEP="TRUE" *) wire n6202_o;
  (* KEEP="TRUE" *) wire n6204_o;
  (* KEEP="TRUE" *) wire n6205_o;
  (* KEEP="TRUE" *) wire n6206_o;
  (* KEEP="TRUE" *) wire n6208_o;
  (* KEEP="TRUE" *) wire n6212_o;
  (* KEEP="TRUE" *) wire n6213_o;
  (* KEEP="TRUE" *) wire n6215_o;
  (* KEEP="TRUE" *) wire n6216_o;
  (* KEEP="TRUE" *) wire n6217_o;
  (* KEEP="TRUE" *) wire n6219_o;
  (* KEEP="TRUE" *) wire n6220_o;
  (* KEEP="TRUE" *) wire n6222_o;
  (* KEEP="TRUE" *) wire n6223_o;
  (* KEEP="TRUE" *) wire n6224_o;
  (* KEEP="TRUE" *) wire n6226_o;
  (* KEEP="TRUE" *) wire n6230_o;
  (* KEEP="TRUE" *) wire n6231_o;
  (* KEEP="TRUE" *) wire n6233_o;
  (* KEEP="TRUE" *) wire n6234_o;
  (* KEEP="TRUE" *) wire n6235_o;
  (* KEEP="TRUE" *) wire n6237_o;
  (* KEEP="TRUE" *) wire n6238_o;
  (* KEEP="TRUE" *) wire n6240_o;
  (* KEEP="TRUE" *) wire n6241_o;
  (* KEEP="TRUE" *) wire n6242_o;
  (* KEEP="TRUE" *) wire n6244_o;
  (* KEEP="TRUE" *) wire n6248_o;
  (* KEEP="TRUE" *) wire n6249_o;
  (* KEEP="TRUE" *) wire n6251_o;
  (* KEEP="TRUE" *) wire n6252_o;
  (* KEEP="TRUE" *) wire n6253_o;
  (* KEEP="TRUE" *) wire n6255_o;
  (* KEEP="TRUE" *) wire n6256_o;
  (* KEEP="TRUE" *) wire n6258_o;
  (* KEEP="TRUE" *) wire n6259_o;
  (* KEEP="TRUE" *) wire n6260_o;
  (* KEEP="TRUE" *) wire n6262_o;
  (* KEEP="TRUE" *) wire n6266_o;
  (* KEEP="TRUE" *) wire n6267_o;
  (* KEEP="TRUE" *) wire n6269_o;
  (* KEEP="TRUE" *) wire n6270_o;
  (* KEEP="TRUE" *) wire n6271_o;
  (* KEEP="TRUE" *) wire n6273_o;
  (* KEEP="TRUE" *) wire n6274_o;
  (* KEEP="TRUE" *) wire n6276_o;
  (* KEEP="TRUE" *) wire n6277_o;
  (* KEEP="TRUE" *) wire n6278_o;
  (* KEEP="TRUE" *) wire n6280_o;
  (* KEEP="TRUE" *) wire n6284_o;
  (* KEEP="TRUE" *) wire n6285_o;
  (* KEEP="TRUE" *) wire n6287_o;
  (* KEEP="TRUE" *) wire n6288_o;
  (* KEEP="TRUE" *) wire n6289_o;
  (* KEEP="TRUE" *) wire n6291_o;
  (* KEEP="TRUE" *) wire n6292_o;
  (* KEEP="TRUE" *) wire n6294_o;
  (* KEEP="TRUE" *) wire n6295_o;
  (* KEEP="TRUE" *) wire n6296_o;
  (* KEEP="TRUE" *) wire n6298_o;
  (* KEEP="TRUE" *) wire n6302_o;
  (* KEEP="TRUE" *) wire n6303_o;
  (* KEEP="TRUE" *) wire n6305_o;
  (* KEEP="TRUE" *) wire n6306_o;
  (* KEEP="TRUE" *) wire n6307_o;
  (* KEEP="TRUE" *) wire n6309_o;
  (* KEEP="TRUE" *) wire n6310_o;
  (* KEEP="TRUE" *) wire n6312_o;
  (* KEEP="TRUE" *) wire n6313_o;
  (* KEEP="TRUE" *) wire n6314_o;
  (* KEEP="TRUE" *) wire n6316_o;
  (* KEEP="TRUE" *) wire n6320_o;
  (* KEEP="TRUE" *) wire n6321_o;
  (* KEEP="TRUE" *) wire n6323_o;
  (* KEEP="TRUE" *) wire n6324_o;
  (* KEEP="TRUE" *) wire n6325_o;
  (* KEEP="TRUE" *) wire n6327_o;
  (* KEEP="TRUE" *) wire n6328_o;
  (* KEEP="TRUE" *) wire n6330_o;
  (* KEEP="TRUE" *) wire n6331_o;
  (* KEEP="TRUE" *) wire n6332_o;
  (* KEEP="TRUE" *) wire n6334_o;
  (* KEEP="TRUE" *) wire n6338_o;
  (* KEEP="TRUE" *) wire n6339_o;
  (* KEEP="TRUE" *) wire n6341_o;
  (* KEEP="TRUE" *) wire n6342_o;
  (* KEEP="TRUE" *) wire n6343_o;
  (* KEEP="TRUE" *) wire n6345_o;
  (* KEEP="TRUE" *) wire n6346_o;
  (* KEEP="TRUE" *) wire n6348_o;
  (* KEEP="TRUE" *) wire n6349_o;
  (* KEEP="TRUE" *) wire n6350_o;
  (* KEEP="TRUE" *) wire n6352_o;
  (* KEEP="TRUE" *) wire n6356_o;
  (* KEEP="TRUE" *) wire n6357_o;
  (* KEEP="TRUE" *) wire n6359_o;
  (* KEEP="TRUE" *) wire n6360_o;
  (* KEEP="TRUE" *) wire n6361_o;
  (* KEEP="TRUE" *) wire n6363_o;
  (* KEEP="TRUE" *) wire n6364_o;
  (* KEEP="TRUE" *) wire n6366_o;
  (* KEEP="TRUE" *) wire n6367_o;
  (* KEEP="TRUE" *) wire n6368_o;
  (* KEEP="TRUE" *) wire n6370_o;
  (* KEEP="TRUE" *) wire n6374_o;
  (* KEEP="TRUE" *) wire n6375_o;
  (* KEEP="TRUE" *) wire n6377_o;
  (* KEEP="TRUE" *) wire n6378_o;
  (* KEEP="TRUE" *) wire n6379_o;
  (* KEEP="TRUE" *) wire n6381_o;
  (* KEEP="TRUE" *) wire n6382_o;
  (* KEEP="TRUE" *) wire n6384_o;
  (* KEEP="TRUE" *) wire n6385_o;
  (* KEEP="TRUE" *) wire n6386_o;
  (* KEEP="TRUE" *) wire n6388_o;
  (* KEEP="TRUE" *) wire n6392_o;
  (* KEEP="TRUE" *) wire n6393_o;
  (* KEEP="TRUE" *) wire n6395_o;
  (* KEEP="TRUE" *) wire n6396_o;
  (* KEEP="TRUE" *) wire n6397_o;
  (* KEEP="TRUE" *) wire n6399_o;
  (* KEEP="TRUE" *) wire n6400_o;
  (* KEEP="TRUE" *) wire n6402_o;
  (* KEEP="TRUE" *) wire n6403_o;
  (* KEEP="TRUE" *) wire n6404_o;
  (* KEEP="TRUE" *) wire n6406_o;
  (* KEEP="TRUE" *) wire n6410_o;
  (* KEEP="TRUE" *) wire n6411_o;
  (* KEEP="TRUE" *) wire n6413_o;
  (* KEEP="TRUE" *) wire n6414_o;
  (* KEEP="TRUE" *) wire n6415_o;
  (* KEEP="TRUE" *) wire n6417_o;
  (* KEEP="TRUE" *) wire n6418_o;
  (* KEEP="TRUE" *) wire n6420_o;
  (* KEEP="TRUE" *) wire n6421_o;
  (* KEEP="TRUE" *) wire n6422_o;
  (* KEEP="TRUE" *) wire n6424_o;
  (* KEEP="TRUE" *) wire n6428_o;
  (* KEEP="TRUE" *) wire n6429_o;
  (* KEEP="TRUE" *) wire n6431_o;
  (* KEEP="TRUE" *) wire n6432_o;
  (* KEEP="TRUE" *) wire n6433_o;
  (* KEEP="TRUE" *) wire n6435_o;
  (* KEEP="TRUE" *) wire n6436_o;
  (* KEEP="TRUE" *) wire n6438_o;
  (* KEEP="TRUE" *) wire n6439_o;
  (* KEEP="TRUE" *) wire n6440_o;
  (* KEEP="TRUE" *) wire n6442_o;
  (* KEEP="TRUE" *) wire n6446_o;
  (* KEEP="TRUE" *) wire n6447_o;
  (* KEEP="TRUE" *) wire n6449_o;
  (* KEEP="TRUE" *) wire n6450_o;
  (* KEEP="TRUE" *) wire n6451_o;
  (* KEEP="TRUE" *) wire n6453_o;
  (* KEEP="TRUE" *) wire n6454_o;
  (* KEEP="TRUE" *) wire n6456_o;
  (* KEEP="TRUE" *) wire n6457_o;
  (* KEEP="TRUE" *) wire n6458_o;
  (* KEEP="TRUE" *) wire n6460_o;
  (* KEEP="TRUE" *) wire n6464_o;
  (* KEEP="TRUE" *) wire n6465_o;
  (* KEEP="TRUE" *) wire n6467_o;
  (* KEEP="TRUE" *) wire n6468_o;
  (* KEEP="TRUE" *) wire n6469_o;
  (* KEEP="TRUE" *) wire n6471_o;
  (* KEEP="TRUE" *) wire n6472_o;
  (* KEEP="TRUE" *) wire n6474_o;
  (* KEEP="TRUE" *) wire n6475_o;
  (* KEEP="TRUE" *) wire n6476_o;
  (* KEEP="TRUE" *) wire n6478_o;
  (* KEEP="TRUE" *) wire n6482_o;
  (* KEEP="TRUE" *) wire n6483_o;
  (* KEEP="TRUE" *) wire n6485_o;
  (* KEEP="TRUE" *) wire n6486_o;
  (* KEEP="TRUE" *) wire n6487_o;
  (* KEEP="TRUE" *) wire n6489_o;
  (* KEEP="TRUE" *) wire n6490_o;
  (* KEEP="TRUE" *) wire n6492_o;
  (* KEEP="TRUE" *) wire n6493_o;
  (* KEEP="TRUE" *) wire n6494_o;
  (* KEEP="TRUE" *) wire n6496_o;
  (* KEEP="TRUE" *) wire n6500_o;
  (* KEEP="TRUE" *) wire n6501_o;
  (* KEEP="TRUE" *) wire n6503_o;
  (* KEEP="TRUE" *) wire n6504_o;
  (* KEEP="TRUE" *) wire n6505_o;
  (* KEEP="TRUE" *) wire n6507_o;
  (* KEEP="TRUE" *) wire n6508_o;
  (* KEEP="TRUE" *) wire n6510_o;
  (* KEEP="TRUE" *) wire n6511_o;
  (* KEEP="TRUE" *) wire n6512_o;
  (* KEEP="TRUE" *) wire n6514_o;
  (* KEEP="TRUE" *) wire n6518_o;
  (* KEEP="TRUE" *) wire n6519_o;
  (* KEEP="TRUE" *) wire n6521_o;
  (* KEEP="TRUE" *) wire n6522_o;
  (* KEEP="TRUE" *) wire n6523_o;
  (* KEEP="TRUE" *) wire n6525_o;
  (* KEEP="TRUE" *) wire n6526_o;
  (* KEEP="TRUE" *) wire n6528_o;
  (* KEEP="TRUE" *) wire n6529_o;
  (* KEEP="TRUE" *) wire n6530_o;
  (* KEEP="TRUE" *) wire n6532_o;
  (* KEEP="TRUE" *) wire n6536_o;
  (* KEEP="TRUE" *) wire n6537_o;
  (* KEEP="TRUE" *) wire n6539_o;
  (* KEEP="TRUE" *) wire n6540_o;
  (* KEEP="TRUE" *) wire n6541_o;
  (* KEEP="TRUE" *) wire n6543_o;
  (* KEEP="TRUE" *) wire n6544_o;
  (* KEEP="TRUE" *) wire n6546_o;
  (* KEEP="TRUE" *) wire n6547_o;
  (* KEEP="TRUE" *) wire n6548_o;
  (* KEEP="TRUE" *) wire n6550_o;
  (* KEEP="TRUE" *) wire n6554_o;
  (* KEEP="TRUE" *) wire n6555_o;
  (* KEEP="TRUE" *) wire n6557_o;
  (* KEEP="TRUE" *) wire n6558_o;
  (* KEEP="TRUE" *) wire n6559_o;
  (* KEEP="TRUE" *) wire n6561_o;
  (* KEEP="TRUE" *) wire n6562_o;
  (* KEEP="TRUE" *) wire n6564_o;
  (* KEEP="TRUE" *) wire n6565_o;
  (* KEEP="TRUE" *) wire n6566_o;
  (* KEEP="TRUE" *) wire n6568_o;
  (* KEEP="TRUE" *) wire n6572_o;
  (* KEEP="TRUE" *) wire n6573_o;
  (* KEEP="TRUE" *) wire n6575_o;
  (* KEEP="TRUE" *) wire n6576_o;
  (* KEEP="TRUE" *) wire n6577_o;
  (* KEEP="TRUE" *) wire n6579_o;
  (* KEEP="TRUE" *) wire n6580_o;
  (* KEEP="TRUE" *) wire n6582_o;
  (* KEEP="TRUE" *) wire n6583_o;
  (* KEEP="TRUE" *) wire n6584_o;
  (* KEEP="TRUE" *) wire n6586_o;
  (* KEEP="TRUE" *) wire n6590_o;
  (* KEEP="TRUE" *) wire n6591_o;
  (* KEEP="TRUE" *) wire n6593_o;
  (* KEEP="TRUE" *) wire n6594_o;
  (* KEEP="TRUE" *) wire n6595_o;
  (* KEEP="TRUE" *) wire n6597_o;
  (* KEEP="TRUE" *) wire n6598_o;
  (* KEEP="TRUE" *) wire n6600_o;
  (* KEEP="TRUE" *) wire n6601_o;
  (* KEEP="TRUE" *) wire n6602_o;
  (* KEEP="TRUE" *) wire n6604_o;
  (* KEEP="TRUE" *) wire n6608_o;
  (* KEEP="TRUE" *) wire n6609_o;
  (* KEEP="TRUE" *) wire n6611_o;
  (* KEEP="TRUE" *) wire n6612_o;
  (* KEEP="TRUE" *) wire n6613_o;
  (* KEEP="TRUE" *) wire n6615_o;
  (* KEEP="TRUE" *) wire n6616_o;
  (* KEEP="TRUE" *) wire n6618_o;
  (* KEEP="TRUE" *) wire n6619_o;
  (* KEEP="TRUE" *) wire n6620_o;
  (* KEEP="TRUE" *) wire n6622_o;
  (* KEEP="TRUE" *) wire n6626_o;
  (* KEEP="TRUE" *) wire n6627_o;
  (* KEEP="TRUE" *) wire n6629_o;
  (* KEEP="TRUE" *) wire n6630_o;
  (* KEEP="TRUE" *) wire n6631_o;
  (* KEEP="TRUE" *) wire n6633_o;
  (* KEEP="TRUE" *) wire n6634_o;
  (* KEEP="TRUE" *) wire n6636_o;
  (* KEEP="TRUE" *) wire n6637_o;
  (* KEEP="TRUE" *) wire n6638_o;
  (* KEEP="TRUE" *) wire n6640_o;
  (* KEEP="TRUE" *) wire n6644_o;
  (* KEEP="TRUE" *) wire n6645_o;
  (* KEEP="TRUE" *) wire n6647_o;
  (* KEEP="TRUE" *) wire n6648_o;
  (* KEEP="TRUE" *) wire n6649_o;
  (* KEEP="TRUE" *) wire n6651_o;
  (* KEEP="TRUE" *) wire n6652_o;
  (* KEEP="TRUE" *) wire n6654_o;
  (* KEEP="TRUE" *) wire n6655_o;
  (* KEEP="TRUE" *) wire n6656_o;
  (* KEEP="TRUE" *) wire n6658_o;
  (* KEEP="TRUE" *) wire n6662_o;
  (* KEEP="TRUE" *) wire n6663_o;
  (* KEEP="TRUE" *) wire n6665_o;
  (* KEEP="TRUE" *) wire n6666_o;
  (* KEEP="TRUE" *) wire n6667_o;
  (* KEEP="TRUE" *) wire n6669_o;
  (* KEEP="TRUE" *) wire n6670_o;
  (* KEEP="TRUE" *) wire n6672_o;
  (* KEEP="TRUE" *) wire n6673_o;
  (* KEEP="TRUE" *) wire n6674_o;
  (* KEEP="TRUE" *) wire n6676_o;
  (* KEEP="TRUE" *) wire n6680_o;
  (* KEEP="TRUE" *) wire n6681_o;
  (* KEEP="TRUE" *) wire n6683_o;
  (* KEEP="TRUE" *) wire n6684_o;
  (* KEEP="TRUE" *) wire n6685_o;
  (* KEEP="TRUE" *) wire n6687_o;
  (* KEEP="TRUE" *) wire n6688_o;
  (* KEEP="TRUE" *) wire n6690_o;
  (* KEEP="TRUE" *) wire n6691_o;
  (* KEEP="TRUE" *) wire n6692_o;
  (* KEEP="TRUE" *) wire n6694_o;
  (* KEEP="TRUE" *) wire n6698_o;
  (* KEEP="TRUE" *) wire n6699_o;
  (* KEEP="TRUE" *) wire n6701_o;
  (* KEEP="TRUE" *) wire n6702_o;
  (* KEEP="TRUE" *) wire n6703_o;
  (* KEEP="TRUE" *) wire n6705_o;
  (* KEEP="TRUE" *) wire n6706_o;
  (* KEEP="TRUE" *) wire n6708_o;
  (* KEEP="TRUE" *) wire n6709_o;
  (* KEEP="TRUE" *) wire n6710_o;
  (* KEEP="TRUE" *) wire n6712_o;
  (* KEEP="TRUE" *) wire n6716_o;
  (* KEEP="TRUE" *) wire n6717_o;
  (* KEEP="TRUE" *) wire n6719_o;
  (* KEEP="TRUE" *) wire n6720_o;
  (* KEEP="TRUE" *) wire n6721_o;
  (* KEEP="TRUE" *) wire n6723_o;
  (* KEEP="TRUE" *) wire n6724_o;
  (* KEEP="TRUE" *) wire n6726_o;
  (* KEEP="TRUE" *) wire n6727_o;
  (* KEEP="TRUE" *) wire n6728_o;
  (* KEEP="TRUE" *) wire n6730_o;
  (* KEEP="TRUE" *) wire n6734_o;
  (* KEEP="TRUE" *) wire n6735_o;
  (* KEEP="TRUE" *) wire n6737_o;
  (* KEEP="TRUE" *) wire n6738_o;
  (* KEEP="TRUE" *) wire n6739_o;
  (* KEEP="TRUE" *) wire n6741_o;
  (* KEEP="TRUE" *) wire n6742_o;
  (* KEEP="TRUE" *) wire n6744_o;
  (* KEEP="TRUE" *) wire n6745_o;
  (* KEEP="TRUE" *) wire n6746_o;
  (* KEEP="TRUE" *) wire n6748_o;
  (* KEEP="TRUE" *) wire n6752_o;
  (* KEEP="TRUE" *) wire n6753_o;
  (* KEEP="TRUE" *) wire n6755_o;
  (* KEEP="TRUE" *) wire n6756_o;
  (* KEEP="TRUE" *) wire n6757_o;
  (* KEEP="TRUE" *) wire n6759_o;
  (* KEEP="TRUE" *) wire n6760_o;
  (* KEEP="TRUE" *) wire n6762_o;
  (* KEEP="TRUE" *) wire n6763_o;
  (* KEEP="TRUE" *) wire n6764_o;
  (* KEEP="TRUE" *) wire n6766_o;
  (* KEEP="TRUE" *) wire n6770_o;
  (* KEEP="TRUE" *) wire n6771_o;
  (* KEEP="TRUE" *) wire n6773_o;
  (* KEEP="TRUE" *) wire n6774_o;
  (* KEEP="TRUE" *) wire n6775_o;
  (* KEEP="TRUE" *) wire n6777_o;
  (* KEEP="TRUE" *) wire n6778_o;
  (* KEEP="TRUE" *) wire n6780_o;
  (* KEEP="TRUE" *) wire n6781_o;
  (* KEEP="TRUE" *) wire n6782_o;
  (* KEEP="TRUE" *) wire n6784_o;
  (* KEEP="TRUE" *) wire n6788_o;
  (* KEEP="TRUE" *) wire n6789_o;
  (* KEEP="TRUE" *) wire n6791_o;
  (* KEEP="TRUE" *) wire n6792_o;
  (* KEEP="TRUE" *) wire n6793_o;
  (* KEEP="TRUE" *) wire n6795_o;
  (* KEEP="TRUE" *) wire n6796_o;
  (* KEEP="TRUE" *) wire n6798_o;
  (* KEEP="TRUE" *) wire n6799_o;
  (* KEEP="TRUE" *) wire n6800_o;
  (* KEEP="TRUE" *) wire n6802_o;
  (* KEEP="TRUE" *) wire n6806_o;
  (* KEEP="TRUE" *) wire n6807_o;
  (* KEEP="TRUE" *) wire n6809_o;
  (* KEEP="TRUE" *) wire n6810_o;
  (* KEEP="TRUE" *) wire n6811_o;
  (* KEEP="TRUE" *) wire n6813_o;
  (* KEEP="TRUE" *) wire n6814_o;
  (* KEEP="TRUE" *) wire n6816_o;
  (* KEEP="TRUE" *) wire n6817_o;
  (* KEEP="TRUE" *) wire n6818_o;
  (* KEEP="TRUE" *) wire n6820_o;
  (* KEEP="TRUE" *) wire n6824_o;
  (* KEEP="TRUE" *) wire n6825_o;
  (* KEEP="TRUE" *) wire n6827_o;
  (* KEEP="TRUE" *) wire n6828_o;
  (* KEEP="TRUE" *) wire n6829_o;
  (* KEEP="TRUE" *) wire n6831_o;
  (* KEEP="TRUE" *) wire n6832_o;
  (* KEEP="TRUE" *) wire n6834_o;
  (* KEEP="TRUE" *) wire n6835_o;
  (* KEEP="TRUE" *) wire n6836_o;
  (* KEEP="TRUE" *) wire n6838_o;
  (* KEEP="TRUE" *) wire n6842_o;
  (* KEEP="TRUE" *) wire n6843_o;
  (* KEEP="TRUE" *) wire n6845_o;
  (* KEEP="TRUE" *) wire n6846_o;
  (* KEEP="TRUE" *) wire n6847_o;
  (* KEEP="TRUE" *) wire n6849_o;
  (* KEEP="TRUE" *) wire n6850_o;
  (* KEEP="TRUE" *) wire n6852_o;
  (* KEEP="TRUE" *) wire n6853_o;
  (* KEEP="TRUE" *) wire n6854_o;
  (* KEEP="TRUE" *) wire n6856_o;
  (* KEEP="TRUE" *) wire n6860_o;
  (* KEEP="TRUE" *) wire n6861_o;
  (* KEEP="TRUE" *) wire n6863_o;
  (* KEEP="TRUE" *) wire n6864_o;
  (* KEEP="TRUE" *) wire n6865_o;
  (* KEEP="TRUE" *) wire n6867_o;
  (* KEEP="TRUE" *) wire n6868_o;
  (* KEEP="TRUE" *) wire n6870_o;
  (* KEEP="TRUE" *) wire n6871_o;
  (* KEEP="TRUE" *) wire n6872_o;
  (* KEEP="TRUE" *) wire n6874_o;
  (* KEEP="TRUE" *) wire n6878_o;
  (* KEEP="TRUE" *) wire n6879_o;
  (* KEEP="TRUE" *) wire n6881_o;
  (* KEEP="TRUE" *) wire n6882_o;
  (* KEEP="TRUE" *) wire n6883_o;
  (* KEEP="TRUE" *) wire n6885_o;
  (* KEEP="TRUE" *) wire n6886_o;
  (* KEEP="TRUE" *) wire n6888_o;
  (* KEEP="TRUE" *) wire n6889_o;
  (* KEEP="TRUE" *) wire n6890_o;
  (* KEEP="TRUE" *) wire n6892_o;
  (* KEEP="TRUE" *) wire n6896_o;
  (* KEEP="TRUE" *) wire n6897_o;
  (* KEEP="TRUE" *) wire n6899_o;
  (* KEEP="TRUE" *) wire n6900_o;
  (* KEEP="TRUE" *) wire n6901_o;
  (* KEEP="TRUE" *) wire n6903_o;
  (* KEEP="TRUE" *) wire n6904_o;
  (* KEEP="TRUE" *) wire n6906_o;
  (* KEEP="TRUE" *) wire n6907_o;
  (* KEEP="TRUE" *) wire n6908_o;
  (* KEEP="TRUE" *) wire n6910_o;
  (* KEEP="TRUE" *) wire n6914_o;
  (* KEEP="TRUE" *) wire n6915_o;
  (* KEEP="TRUE" *) wire n6917_o;
  (* KEEP="TRUE" *) wire n6918_o;
  (* KEEP="TRUE" *) wire n6919_o;
  (* KEEP="TRUE" *) wire n6921_o;
  (* KEEP="TRUE" *) wire n6922_o;
  (* KEEP="TRUE" *) wire n6924_o;
  (* KEEP="TRUE" *) wire n6925_o;
  (* KEEP="TRUE" *) wire n6926_o;
  (* KEEP="TRUE" *) wire n6928_o;
  (* KEEP="TRUE" *) wire n6932_o;
  (* KEEP="TRUE" *) wire n6933_o;
  (* KEEP="TRUE" *) wire n6935_o;
  (* KEEP="TRUE" *) wire n6936_o;
  (* KEEP="TRUE" *) wire n6937_o;
  (* KEEP="TRUE" *) wire n6939_o;
  (* KEEP="TRUE" *) wire n6940_o;
  (* KEEP="TRUE" *) wire n6942_o;
  (* KEEP="TRUE" *) wire n6943_o;
  (* KEEP="TRUE" *) wire n6944_o;
  (* KEEP="TRUE" *) wire n6946_o;
  (* KEEP="TRUE" *) wire n6950_o;
  (* KEEP="TRUE" *) wire n6951_o;
  (* KEEP="TRUE" *) wire n6953_o;
  (* KEEP="TRUE" *) wire n6954_o;
  (* KEEP="TRUE" *) wire n6955_o;
  (* KEEP="TRUE" *) wire n6957_o;
  (* KEEP="TRUE" *) wire n6958_o;
  (* KEEP="TRUE" *) wire n6960_o;
  (* KEEP="TRUE" *) wire n6961_o;
  (* KEEP="TRUE" *) wire n6962_o;
  (* KEEP="TRUE" *) wire n6964_o;
  (* KEEP="TRUE" *) wire n6968_o;
  (* KEEP="TRUE" *) wire n6969_o;
  (* KEEP="TRUE" *) wire n6971_o;
  (* KEEP="TRUE" *) wire n6972_o;
  (* KEEP="TRUE" *) wire n6973_o;
  (* KEEP="TRUE" *) wire n6975_o;
  (* KEEP="TRUE" *) wire n6976_o;
  (* KEEP="TRUE" *) wire n6978_o;
  (* KEEP="TRUE" *) wire n6979_o;
  (* KEEP="TRUE" *) wire n6980_o;
  (* KEEP="TRUE" *) wire n6982_o;
  (* KEEP="TRUE" *) wire n6986_o;
  (* KEEP="TRUE" *) wire n6987_o;
  (* KEEP="TRUE" *) wire n6989_o;
  (* KEEP="TRUE" *) wire n6990_o;
  (* KEEP="TRUE" *) wire n6991_o;
  (* KEEP="TRUE" *) wire n6993_o;
  (* KEEP="TRUE" *) wire n6994_o;
  (* KEEP="TRUE" *) wire n6996_o;
  (* KEEP="TRUE" *) wire n6997_o;
  (* KEEP="TRUE" *) wire n6998_o;
  (* KEEP="TRUE" *) wire n7000_o;
  (* KEEP="TRUE" *) wire n7004_o;
  (* KEEP="TRUE" *) wire n7005_o;
  (* KEEP="TRUE" *) wire n7007_o;
  (* KEEP="TRUE" *) wire n7008_o;
  (* KEEP="TRUE" *) wire n7009_o;
  (* KEEP="TRUE" *) wire n7011_o;
  (* KEEP="TRUE" *) wire n7012_o;
  (* KEEP="TRUE" *) wire n7014_o;
  (* KEEP="TRUE" *) wire n7015_o;
  (* KEEP="TRUE" *) wire n7016_o;
  (* KEEP="TRUE" *) wire n7018_o;
  (* KEEP="TRUE" *) wire n7022_o;
  (* KEEP="TRUE" *) wire n7023_o;
  (* KEEP="TRUE" *) wire n7025_o;
  (* KEEP="TRUE" *) wire n7026_o;
  (* KEEP="TRUE" *) wire n7027_o;
  (* KEEP="TRUE" *) wire n7029_o;
  (* KEEP="TRUE" *) wire n7030_o;
  (* KEEP="TRUE" *) wire n7032_o;
  (* KEEP="TRUE" *) wire n7033_o;
  (* KEEP="TRUE" *) wire n7034_o;
  (* KEEP="TRUE" *) wire n7036_o;
  (* KEEP="TRUE" *) wire n7040_o;
  (* KEEP="TRUE" *) wire n7041_o;
  (* KEEP="TRUE" *) wire n7043_o;
  (* KEEP="TRUE" *) wire n7044_o;
  (* KEEP="TRUE" *) wire n7045_o;
  (* KEEP="TRUE" *) wire n7047_o;
  (* KEEP="TRUE" *) wire n7048_o;
  (* KEEP="TRUE" *) wire n7050_o;
  (* KEEP="TRUE" *) wire n7051_o;
  (* KEEP="TRUE" *) wire n7052_o;
  (* KEEP="TRUE" *) wire n7054_o;
  (* KEEP="TRUE" *) wire n7058_o;
  (* KEEP="TRUE" *) wire n7059_o;
  (* KEEP="TRUE" *) wire n7061_o;
  (* KEEP="TRUE" *) wire n7062_o;
  (* KEEP="TRUE" *) wire n7063_o;
  (* KEEP="TRUE" *) wire n7065_o;
  (* KEEP="TRUE" *) wire n7066_o;
  (* KEEP="TRUE" *) wire n7068_o;
  (* KEEP="TRUE" *) wire n7069_o;
  (* KEEP="TRUE" *) wire n7070_o;
  (* KEEP="TRUE" *) wire n7072_o;
  (* KEEP="TRUE" *) wire n7076_o;
  (* KEEP="TRUE" *) wire n7077_o;
  (* KEEP="TRUE" *) wire n7079_o;
  (* KEEP="TRUE" *) wire n7080_o;
  (* KEEP="TRUE" *) wire n7081_o;
  (* KEEP="TRUE" *) wire n7083_o;
  (* KEEP="TRUE" *) wire n7084_o;
  (* KEEP="TRUE" *) wire n7086_o;
  (* KEEP="TRUE" *) wire n7087_o;
  (* KEEP="TRUE" *) wire n7088_o;
  (* KEEP="TRUE" *) wire n7090_o;
  (* KEEP="TRUE" *) wire n7094_o;
  (* KEEP="TRUE" *) wire n7095_o;
  (* KEEP="TRUE" *) wire n7097_o;
  (* KEEP="TRUE" *) wire n7098_o;
  (* KEEP="TRUE" *) wire n7099_o;
  (* KEEP="TRUE" *) wire n7101_o;
  (* KEEP="TRUE" *) wire n7102_o;
  (* KEEP="TRUE" *) wire n7104_o;
  (* KEEP="TRUE" *) wire n7105_o;
  (* KEEP="TRUE" *) wire n7106_o;
  (* KEEP="TRUE" *) wire n7108_o;
  (* KEEP="TRUE" *) wire n7112_o;
  (* KEEP="TRUE" *) wire n7113_o;
  (* KEEP="TRUE" *) wire n7115_o;
  (* KEEP="TRUE" *) wire n7116_o;
  (* KEEP="TRUE" *) wire n7117_o;
  (* KEEP="TRUE" *) wire n7119_o;
  (* KEEP="TRUE" *) wire n7120_o;
  (* KEEP="TRUE" *) wire n7122_o;
  (* KEEP="TRUE" *) wire n7123_o;
  (* KEEP="TRUE" *) wire n7124_o;
  (* KEEP="TRUE" *) wire n7126_o;
  (* KEEP="TRUE" *) wire n7130_o;
  (* KEEP="TRUE" *) wire n7131_o;
  (* KEEP="TRUE" *) wire n7133_o;
  (* KEEP="TRUE" *) wire n7134_o;
  (* KEEP="TRUE" *) wire n7135_o;
  (* KEEP="TRUE" *) wire n7137_o;
  (* KEEP="TRUE" *) wire n7138_o;
  (* KEEP="TRUE" *) wire n7140_o;
  (* KEEP="TRUE" *) wire n7141_o;
  (* KEEP="TRUE" *) wire n7142_o;
  (* KEEP="TRUE" *) wire n7144_o;
  (* KEEP="TRUE" *) wire n7148_o;
  (* KEEP="TRUE" *) wire n7149_o;
  (* KEEP="TRUE" *) wire n7151_o;
  (* KEEP="TRUE" *) wire n7152_o;
  (* KEEP="TRUE" *) wire n7153_o;
  (* KEEP="TRUE" *) wire n7155_o;
  (* KEEP="TRUE" *) wire n7156_o;
  (* KEEP="TRUE" *) wire n7158_o;
  (* KEEP="TRUE" *) wire n7159_o;
  (* KEEP="TRUE" *) wire n7160_o;
  (* KEEP="TRUE" *) wire n7162_o;
  (* KEEP="TRUE" *) wire n7166_o;
  (* KEEP="TRUE" *) wire n7167_o;
  (* KEEP="TRUE" *) wire n7169_o;
  (* KEEP="TRUE" *) wire n7170_o;
  (* KEEP="TRUE" *) wire n7171_o;
  (* KEEP="TRUE" *) wire n7173_o;
  (* KEEP="TRUE" *) wire n7174_o;
  (* KEEP="TRUE" *) wire n7176_o;
  (* KEEP="TRUE" *) wire n7177_o;
  (* KEEP="TRUE" *) wire n7178_o;
  (* KEEP="TRUE" *) wire n7180_o;
  (* KEEP="TRUE" *) wire n7184_o;
  (* KEEP="TRUE" *) wire n7185_o;
  (* KEEP="TRUE" *) wire n7187_o;
  (* KEEP="TRUE" *) wire n7188_o;
  (* KEEP="TRUE" *) wire n7189_o;
  (* KEEP="TRUE" *) wire n7191_o;
  (* KEEP="TRUE" *) wire n7192_o;
  (* KEEP="TRUE" *) wire n7194_o;
  (* KEEP="TRUE" *) wire n7195_o;
  (* KEEP="TRUE" *) wire n7196_o;
  (* KEEP="TRUE" *) wire n7198_o;
  (* KEEP="TRUE" *) wire n7202_o;
  (* KEEP="TRUE" *) wire n7203_o;
  (* KEEP="TRUE" *) wire n7205_o;
  (* KEEP="TRUE" *) wire n7206_o;
  (* KEEP="TRUE" *) wire n7207_o;
  (* KEEP="TRUE" *) wire n7209_o;
  (* KEEP="TRUE" *) wire n7210_o;
  (* KEEP="TRUE" *) wire n7212_o;
  (* KEEP="TRUE" *) wire n7213_o;
  (* KEEP="TRUE" *) wire n7214_o;
  (* KEEP="TRUE" *) wire n7216_o;
  (* KEEP="TRUE" *) wire n7220_o;
  (* KEEP="TRUE" *) wire n7221_o;
  (* KEEP="TRUE" *) wire n7223_o;
  (* KEEP="TRUE" *) wire n7224_o;
  (* KEEP="TRUE" *) wire n7225_o;
  (* KEEP="TRUE" *) wire n7227_o;
  (* KEEP="TRUE" *) wire n7228_o;
  (* KEEP="TRUE" *) wire n7230_o;
  (* KEEP="TRUE" *) wire n7231_o;
  (* KEEP="TRUE" *) wire n7232_o;
  (* KEEP="TRUE" *) wire n7234_o;
  (* KEEP="TRUE" *) wire n7238_o;
  (* KEEP="TRUE" *) wire n7239_o;
  (* KEEP="TRUE" *) wire n7241_o;
  (* KEEP="TRUE" *) wire n7242_o;
  (* KEEP="TRUE" *) wire n7243_o;
  (* KEEP="TRUE" *) wire n7245_o;
  (* KEEP="TRUE" *) wire n7246_o;
  (* KEEP="TRUE" *) wire n7248_o;
  (* KEEP="TRUE" *) wire n7249_o;
  (* KEEP="TRUE" *) wire n7250_o;
  (* KEEP="TRUE" *) wire n7252_o;
  (* KEEP="TRUE" *) wire n7256_o;
  (* KEEP="TRUE" *) wire n7257_o;
  (* KEEP="TRUE" *) wire n7259_o;
  (* KEEP="TRUE" *) wire n7260_o;
  (* KEEP="TRUE" *) wire n7261_o;
  (* KEEP="TRUE" *) wire n7263_o;
  (* KEEP="TRUE" *) wire n7264_o;
  (* KEEP="TRUE" *) wire n7266_o;
  (* KEEP="TRUE" *) wire n7267_o;
  (* KEEP="TRUE" *) wire n7268_o;
  (* KEEP="TRUE" *) wire n7270_o;
  (* KEEP="TRUE" *) wire n7274_o;
  (* KEEP="TRUE" *) wire n7275_o;
  (* KEEP="TRUE" *) wire n7277_o;
  (* KEEP="TRUE" *) wire n7278_o;
  (* KEEP="TRUE" *) wire n7279_o;
  (* KEEP="TRUE" *) wire n7281_o;
  (* KEEP="TRUE" *) wire n7282_o;
  (* KEEP="TRUE" *) wire n7284_o;
  (* KEEP="TRUE" *) wire n7285_o;
  (* KEEP="TRUE" *) wire n7286_o;
  (* KEEP="TRUE" *) wire n7288_o;
  (* KEEP="TRUE" *) wire n7292_o;
  (* KEEP="TRUE" *) wire n7293_o;
  (* KEEP="TRUE" *) wire n7295_o;
  (* KEEP="TRUE" *) wire n7296_o;
  (* KEEP="TRUE" *) wire n7297_o;
  (* KEEP="TRUE" *) wire n7299_o;
  (* KEEP="TRUE" *) wire n7300_o;
  (* KEEP="TRUE" *) wire n7302_o;
  (* KEEP="TRUE" *) wire n7303_o;
  (* KEEP="TRUE" *) wire n7304_o;
  (* KEEP="TRUE" *) wire n7306_o;
  (* KEEP="TRUE" *) wire n7310_o;
  (* KEEP="TRUE" *) wire n7311_o;
  (* KEEP="TRUE" *) wire n7313_o;
  (* KEEP="TRUE" *) wire n7314_o;
  (* KEEP="TRUE" *) wire n7315_o;
  (* KEEP="TRUE" *) wire n7317_o;
  (* KEEP="TRUE" *) wire n7318_o;
  (* KEEP="TRUE" *) wire n7320_o;
  (* KEEP="TRUE" *) wire n7321_o;
  (* KEEP="TRUE" *) wire n7322_o;
  (* KEEP="TRUE" *) wire n7324_o;
  (* KEEP="TRUE" *) wire n7328_o;
  (* KEEP="TRUE" *) wire n7329_o;
  (* KEEP="TRUE" *) wire n7331_o;
  (* KEEP="TRUE" *) wire n7332_o;
  (* KEEP="TRUE" *) wire n7333_o;
  (* KEEP="TRUE" *) wire n7335_o;
  (* KEEP="TRUE" *) wire n7336_o;
  (* KEEP="TRUE" *) wire n7338_o;
  (* KEEP="TRUE" *) wire n7339_o;
  (* KEEP="TRUE" *) wire n7340_o;
  (* KEEP="TRUE" *) wire n7342_o;
  (* KEEP="TRUE" *) wire n7346_o;
  (* KEEP="TRUE" *) wire n7347_o;
  (* KEEP="TRUE" *) wire n7349_o;
  (* KEEP="TRUE" *) wire n7350_o;
  (* KEEP="TRUE" *) wire n7351_o;
  (* KEEP="TRUE" *) wire n7353_o;
  (* KEEP="TRUE" *) wire n7354_o;
  (* KEEP="TRUE" *) wire n7356_o;
  (* KEEP="TRUE" *) wire n7357_o;
  (* KEEP="TRUE" *) wire n7358_o;
  (* KEEP="TRUE" *) wire n7360_o;
  (* KEEP="TRUE" *) wire n7364_o;
  (* KEEP="TRUE" *) wire n7365_o;
  (* KEEP="TRUE" *) wire n7367_o;
  (* KEEP="TRUE" *) wire n7368_o;
  (* KEEP="TRUE" *) wire n7369_o;
  (* KEEP="TRUE" *) wire n7371_o;
  (* KEEP="TRUE" *) wire n7372_o;
  (* KEEP="TRUE" *) wire n7374_o;
  (* KEEP="TRUE" *) wire n7375_o;
  (* KEEP="TRUE" *) wire n7376_o;
  (* KEEP="TRUE" *) wire n7378_o;
  (* KEEP="TRUE" *) wire n7382_o;
  (* KEEP="TRUE" *) wire n7383_o;
  (* KEEP="TRUE" *) wire n7385_o;
  (* KEEP="TRUE" *) wire n7386_o;
  (* KEEP="TRUE" *) wire n7387_o;
  (* KEEP="TRUE" *) wire n7389_o;
  (* KEEP="TRUE" *) wire n7390_o;
  (* KEEP="TRUE" *) wire n7392_o;
  (* KEEP="TRUE" *) wire n7393_o;
  (* KEEP="TRUE" *) wire n7394_o;
  (* KEEP="TRUE" *) wire n7396_o;
  (* KEEP="TRUE" *) wire n7400_o;
  (* KEEP="TRUE" *) wire n7401_o;
  (* KEEP="TRUE" *) wire n7403_o;
  (* KEEP="TRUE" *) wire n7404_o;
  (* KEEP="TRUE" *) wire n7405_o;
  (* KEEP="TRUE" *) wire n7407_o;
  (* KEEP="TRUE" *) wire n7408_o;
  (* KEEP="TRUE" *) wire n7410_o;
  (* KEEP="TRUE" *) wire n7411_o;
  (* KEEP="TRUE" *) wire n7412_o;
  (* KEEP="TRUE" *) wire n7414_o;
  (* KEEP="TRUE" *) wire n7418_o;
  (* KEEP="TRUE" *) wire n7419_o;
  (* KEEP="TRUE" *) wire n7421_o;
  (* KEEP="TRUE" *) wire n7422_o;
  (* KEEP="TRUE" *) wire n7423_o;
  (* KEEP="TRUE" *) wire n7425_o;
  (* KEEP="TRUE" *) wire n7426_o;
  (* KEEP="TRUE" *) wire n7428_o;
  (* KEEP="TRUE" *) wire n7429_o;
  (* KEEP="TRUE" *) wire n7430_o;
  (* KEEP="TRUE" *) wire n7432_o;
  (* KEEP="TRUE" *) wire n7436_o;
  (* KEEP="TRUE" *) wire n7437_o;
  (* KEEP="TRUE" *) wire n7439_o;
  (* KEEP="TRUE" *) wire n7440_o;
  (* KEEP="TRUE" *) wire n7441_o;
  (* KEEP="TRUE" *) wire n7443_o;
  (* KEEP="TRUE" *) wire n7444_o;
  (* KEEP="TRUE" *) wire n7446_o;
  (* KEEP="TRUE" *) wire n7447_o;
  (* KEEP="TRUE" *) wire n7448_o;
  (* KEEP="TRUE" *) wire n7450_o;
  (* KEEP="TRUE" *) wire n7454_o;
  (* KEEP="TRUE" *) wire n7455_o;
  (* KEEP="TRUE" *) wire n7457_o;
  (* KEEP="TRUE" *) wire n7458_o;
  (* KEEP="TRUE" *) wire n7459_o;
  (* KEEP="TRUE" *) wire n7461_o;
  (* KEEP="TRUE" *) wire n7462_o;
  (* KEEP="TRUE" *) wire n7464_o;
  (* KEEP="TRUE" *) wire n7465_o;
  (* KEEP="TRUE" *) wire n7466_o;
  (* KEEP="TRUE" *) wire n7468_o;
  (* KEEP="TRUE" *) wire n7472_o;
  (* KEEP="TRUE" *) wire n7473_o;
  (* KEEP="TRUE" *) wire n7475_o;
  (* KEEP="TRUE" *) wire n7476_o;
  (* KEEP="TRUE" *) wire n7477_o;
  (* KEEP="TRUE" *) wire n7479_o;
  (* KEEP="TRUE" *) wire n7480_o;
  (* KEEP="TRUE" *) wire n7482_o;
  (* KEEP="TRUE" *) wire n7483_o;
  (* KEEP="TRUE" *) wire n7484_o;
  (* KEEP="TRUE" *) wire n7486_o;
  (* KEEP="TRUE" *) wire n7490_o;
  (* KEEP="TRUE" *) wire n7491_o;
  (* KEEP="TRUE" *) wire n7493_o;
  (* KEEP="TRUE" *) wire n7494_o;
  (* KEEP="TRUE" *) wire n7495_o;
  (* KEEP="TRUE" *) wire n7497_o;
  (* KEEP="TRUE" *) wire n7498_o;
  (* KEEP="TRUE" *) wire n7500_o;
  (* KEEP="TRUE" *) wire n7501_o;
  (* KEEP="TRUE" *) wire n7502_o;
  (* KEEP="TRUE" *) wire n7504_o;
  (* KEEP="TRUE" *) wire n7508_o;
  (* KEEP="TRUE" *) wire n7509_o;
  (* KEEP="TRUE" *) wire n7511_o;
  (* KEEP="TRUE" *) wire n7512_o;
  (* KEEP="TRUE" *) wire n7513_o;
  (* KEEP="TRUE" *) wire n7515_o;
  (* KEEP="TRUE" *) wire n7516_o;
  (* KEEP="TRUE" *) wire n7518_o;
  (* KEEP="TRUE" *) wire n7519_o;
  (* KEEP="TRUE" *) wire n7520_o;
  (* KEEP="TRUE" *) wire n7522_o;
  (* KEEP="TRUE" *) wire n7526_o;
  (* KEEP="TRUE" *) wire n7527_o;
  (* KEEP="TRUE" *) wire n7529_o;
  (* KEEP="TRUE" *) wire n7530_o;
  (* KEEP="TRUE" *) wire n7531_o;
  (* KEEP="TRUE" *) wire n7533_o;
  (* KEEP="TRUE" *) wire n7534_o;
  (* KEEP="TRUE" *) wire n7536_o;
  (* KEEP="TRUE" *) wire n7537_o;
  (* KEEP="TRUE" *) wire n7538_o;
  (* KEEP="TRUE" *) wire n7540_o;
  (* KEEP="TRUE" *) wire n7544_o;
  (* KEEP="TRUE" *) wire n7545_o;
  (* KEEP="TRUE" *) wire n7547_o;
  (* KEEP="TRUE" *) wire n7548_o;
  (* KEEP="TRUE" *) wire n7549_o;
  (* KEEP="TRUE" *) wire n7551_o;
  (* KEEP="TRUE" *) wire n7552_o;
  (* KEEP="TRUE" *) wire n7554_o;
  (* KEEP="TRUE" *) wire n7555_o;
  (* KEEP="TRUE" *) wire n7556_o;
  (* KEEP="TRUE" *) wire n7558_o;
  (* KEEP="TRUE" *) wire n7562_o;
  (* KEEP="TRUE" *) wire n7563_o;
  (* KEEP="TRUE" *) wire n7565_o;
  (* KEEP="TRUE" *) wire n7566_o;
  (* KEEP="TRUE" *) wire n7567_o;
  (* KEEP="TRUE" *) wire n7569_o;
  (* KEEP="TRUE" *) wire n7570_o;
  (* KEEP="TRUE" *) wire n7572_o;
  (* KEEP="TRUE" *) wire n7573_o;
  (* KEEP="TRUE" *) wire n7574_o;
  (* KEEP="TRUE" *) wire n7576_o;
  (* KEEP="TRUE" *) wire n7580_o;
  (* KEEP="TRUE" *) wire n7581_o;
  (* KEEP="TRUE" *) wire n7583_o;
  (* KEEP="TRUE" *) wire n7584_o;
  (* KEEP="TRUE" *) wire n7585_o;
  (* KEEP="TRUE" *) wire n7587_o;
  (* KEEP="TRUE" *) wire n7588_o;
  (* KEEP="TRUE" *) wire n7590_o;
  (* KEEP="TRUE" *) wire n7591_o;
  (* KEEP="TRUE" *) wire n7592_o;
  (* KEEP="TRUE" *) wire n7594_o;
  (* KEEP="TRUE" *) wire n7598_o;
  (* KEEP="TRUE" *) wire n7599_o;
  (* KEEP="TRUE" *) wire n7601_o;
  (* KEEP="TRUE" *) wire n7602_o;
  (* KEEP="TRUE" *) wire n7603_o;
  (* KEEP="TRUE" *) wire n7605_o;
  (* KEEP="TRUE" *) wire n7606_o;
  (* KEEP="TRUE" *) wire n7608_o;
  (* KEEP="TRUE" *) wire n7609_o;
  (* KEEP="TRUE" *) wire n7610_o;
  (* KEEP="TRUE" *) wire n7612_o;
  (* KEEP="TRUE" *) wire n7616_o;
  (* KEEP="TRUE" *) wire n7617_o;
  (* KEEP="TRUE" *) wire n7619_o;
  (* KEEP="TRUE" *) wire n7620_o;
  (* KEEP="TRUE" *) wire n7621_o;
  (* KEEP="TRUE" *) wire n7623_o;
  (* KEEP="TRUE" *) wire n7624_o;
  (* KEEP="TRUE" *) wire n7626_o;
  (* KEEP="TRUE" *) wire n7627_o;
  (* KEEP="TRUE" *) wire n7628_o;
  (* KEEP="TRUE" *) wire n7630_o;
  (* KEEP="TRUE" *) wire n7634_o;
  (* KEEP="TRUE" *) wire n7635_o;
  (* KEEP="TRUE" *) wire n7637_o;
  (* KEEP="TRUE" *) wire n7638_o;
  (* KEEP="TRUE" *) wire n7639_o;
  (* KEEP="TRUE" *) wire n7641_o;
  (* KEEP="TRUE" *) wire n7642_o;
  (* KEEP="TRUE" *) wire n7644_o;
  (* KEEP="TRUE" *) wire n7645_o;
  (* KEEP="TRUE" *) wire n7646_o;
  (* KEEP="TRUE" *) wire n7648_o;
  (* KEEP="TRUE" *) wire n7652_o;
  (* KEEP="TRUE" *) wire n7653_o;
  (* KEEP="TRUE" *) wire n7655_o;
  (* KEEP="TRUE" *) wire n7656_o;
  (* KEEP="TRUE" *) wire n7657_o;
  (* KEEP="TRUE" *) wire n7659_o;
  (* KEEP="TRUE" *) wire n7660_o;
  (* KEEP="TRUE" *) wire n7662_o;
  (* KEEP="TRUE" *) wire n7663_o;
  (* KEEP="TRUE" *) wire n7664_o;
  (* KEEP="TRUE" *) wire n7666_o;
  (* KEEP="TRUE" *) wire n7670_o;
  (* KEEP="TRUE" *) wire n7671_o;
  (* KEEP="TRUE" *) wire n7673_o;
  (* KEEP="TRUE" *) wire n7674_o;
  (* KEEP="TRUE" *) wire n7675_o;
  (* KEEP="TRUE" *) wire n7677_o;
  (* KEEP="TRUE" *) wire n7678_o;
  (* KEEP="TRUE" *) wire n7680_o;
  (* KEEP="TRUE" *) wire n7681_o;
  (* KEEP="TRUE" *) wire n7682_o;
  (* KEEP="TRUE" *) wire n7684_o;
  (* KEEP="TRUE" *) wire n7688_o;
  (* KEEP="TRUE" *) wire n7689_o;
  (* KEEP="TRUE" *) wire n7691_o;
  (* KEEP="TRUE" *) wire n7692_o;
  (* KEEP="TRUE" *) wire n7693_o;
  (* KEEP="TRUE" *) wire n7695_o;
  (* KEEP="TRUE" *) wire n7696_o;
  (* KEEP="TRUE" *) wire n7698_o;
  (* KEEP="TRUE" *) wire n7699_o;
  (* KEEP="TRUE" *) wire n7700_o;
  (* KEEP="TRUE" *) wire n7702_o;
  (* KEEP="TRUE" *) wire n7706_o;
  (* KEEP="TRUE" *) wire n7707_o;
  (* KEEP="TRUE" *) wire n7709_o;
  (* KEEP="TRUE" *) wire n7710_o;
  (* KEEP="TRUE" *) wire n7711_o;
  (* KEEP="TRUE" *) wire n7713_o;
  (* KEEP="TRUE" *) wire n7714_o;
  (* KEEP="TRUE" *) wire n7716_o;
  (* KEEP="TRUE" *) wire n7717_o;
  (* KEEP="TRUE" *) wire n7718_o;
  (* KEEP="TRUE" *) wire n7720_o;
  (* KEEP="TRUE" *) wire n7724_o;
  (* KEEP="TRUE" *) wire n7725_o;
  (* KEEP="TRUE" *) wire n7727_o;
  (* KEEP="TRUE" *) wire n7728_o;
  (* KEEP="TRUE" *) wire n7729_o;
  (* KEEP="TRUE" *) wire n7731_o;
  (* KEEP="TRUE" *) wire n7732_o;
  (* KEEP="TRUE" *) wire n7734_o;
  (* KEEP="TRUE" *) wire n7735_o;
  (* KEEP="TRUE" *) wire n7736_o;
  (* KEEP="TRUE" *) wire n7738_o;
  (* KEEP="TRUE" *) wire n7742_o;
  (* KEEP="TRUE" *) wire n7743_o;
  (* KEEP="TRUE" *) wire n7745_o;
  (* KEEP="TRUE" *) wire n7746_o;
  (* KEEP="TRUE" *) wire n7747_o;
  (* KEEP="TRUE" *) wire n7749_o;
  (* KEEP="TRUE" *) wire n7750_o;
  (* KEEP="TRUE" *) wire n7752_o;
  (* KEEP="TRUE" *) wire n7753_o;
  (* KEEP="TRUE" *) wire n7754_o;
  (* KEEP="TRUE" *) wire n7756_o;
  (* KEEP="TRUE" *) wire n7760_o;
  (* KEEP="TRUE" *) wire n7761_o;
  (* KEEP="TRUE" *) wire n7763_o;
  (* KEEP="TRUE" *) wire n7764_o;
  (* KEEP="TRUE" *) wire n7765_o;
  (* KEEP="TRUE" *) wire n7767_o;
  (* KEEP="TRUE" *) wire n7768_o;
  (* KEEP="TRUE" *) wire n7770_o;
  (* KEEP="TRUE" *) wire n7771_o;
  (* KEEP="TRUE" *) wire n7772_o;
  (* KEEP="TRUE" *) wire n7774_o;
  (* KEEP="TRUE" *) wire n7778_o;
  (* KEEP="TRUE" *) wire n7779_o;
  (* KEEP="TRUE" *) wire n7781_o;
  (* KEEP="TRUE" *) wire n7782_o;
  (* KEEP="TRUE" *) wire n7783_o;
  (* KEEP="TRUE" *) wire n7785_o;
  (* KEEP="TRUE" *) wire n7786_o;
  (* KEEP="TRUE" *) wire n7788_o;
  (* KEEP="TRUE" *) wire n7789_o;
  (* KEEP="TRUE" *) wire n7790_o;
  (* KEEP="TRUE" *) wire n7792_o;
  (* KEEP="TRUE" *) wire n7796_o;
  (* KEEP="TRUE" *) wire n7797_o;
  (* KEEP="TRUE" *) wire n7799_o;
  (* KEEP="TRUE" *) wire n7800_o;
  (* KEEP="TRUE" *) wire n7801_o;
  (* KEEP="TRUE" *) wire n7803_o;
  (* KEEP="TRUE" *) wire n7804_o;
  (* KEEP="TRUE" *) wire n7806_o;
  (* KEEP="TRUE" *) wire n7807_o;
  (* KEEP="TRUE" *) wire n7808_o;
  (* KEEP="TRUE" *) wire n7810_o;
  (* KEEP="TRUE" *) wire n7814_o;
  (* KEEP="TRUE" *) wire n7815_o;
  (* KEEP="TRUE" *) wire n7817_o;
  (* KEEP="TRUE" *) wire n7818_o;
  (* KEEP="TRUE" *) wire n7819_o;
  (* KEEP="TRUE" *) wire n7821_o;
  (* KEEP="TRUE" *) wire n7822_o;
  (* KEEP="TRUE" *) wire n7824_o;
  (* KEEP="TRUE" *) wire n7825_o;
  (* KEEP="TRUE" *) wire n7826_o;
  (* KEEP="TRUE" *) wire n7828_o;
  (* KEEP="TRUE" *) wire n7832_o;
  (* KEEP="TRUE" *) wire n7833_o;
  (* KEEP="TRUE" *) wire n7835_o;
  (* KEEP="TRUE" *) wire n7836_o;
  (* KEEP="TRUE" *) wire n7837_o;
  (* KEEP="TRUE" *) wire n7839_o;
  (* KEEP="TRUE" *) wire n7840_o;
  (* KEEP="TRUE" *) wire n7842_o;
  (* KEEP="TRUE" *) wire n7843_o;
  (* KEEP="TRUE" *) wire n7844_o;
  (* KEEP="TRUE" *) wire n7846_o;
  (* KEEP="TRUE" *) wire n7850_o;
  (* KEEP="TRUE" *) wire n7851_o;
  (* KEEP="TRUE" *) wire n7853_o;
  (* KEEP="TRUE" *) wire n7854_o;
  (* KEEP="TRUE" *) wire n7855_o;
  (* KEEP="TRUE" *) wire n7857_o;
  (* KEEP="TRUE" *) wire n7858_o;
  (* KEEP="TRUE" *) wire n7860_o;
  (* KEEP="TRUE" *) wire n7861_o;
  (* KEEP="TRUE" *) wire n7862_o;
  (* KEEP="TRUE" *) wire n7864_o;
  (* KEEP="TRUE" *) wire n7868_o;
  (* KEEP="TRUE" *) wire n7869_o;
  (* KEEP="TRUE" *) wire n7871_o;
  (* KEEP="TRUE" *) wire n7872_o;
  (* KEEP="TRUE" *) wire n7873_o;
  (* KEEP="TRUE" *) wire n7875_o;
  (* KEEP="TRUE" *) wire n7876_o;
  (* KEEP="TRUE" *) wire n7878_o;
  (* KEEP="TRUE" *) wire n7879_o;
  (* KEEP="TRUE" *) wire n7880_o;
  (* KEEP="TRUE" *) wire n7882_o;
  (* KEEP="TRUE" *) wire n7886_o;
  (* KEEP="TRUE" *) wire n7887_o;
  (* KEEP="TRUE" *) wire n7889_o;
  (* KEEP="TRUE" *) wire n7890_o;
  (* KEEP="TRUE" *) wire n7891_o;
  (* KEEP="TRUE" *) wire n7893_o;
  (* KEEP="TRUE" *) wire n7894_o;
  (* KEEP="TRUE" *) wire n7896_o;
  (* KEEP="TRUE" *) wire n7897_o;
  (* KEEP="TRUE" *) wire n7898_o;
  (* KEEP="TRUE" *) wire n7900_o;
  (* KEEP="TRUE" *) wire n7904_o;
  (* KEEP="TRUE" *) wire n7905_o;
  (* KEEP="TRUE" *) wire n7907_o;
  (* KEEP="TRUE" *) wire n7908_o;
  (* KEEP="TRUE" *) wire n7909_o;
  (* KEEP="TRUE" *) wire n7911_o;
  (* KEEP="TRUE" *) wire n7912_o;
  (* KEEP="TRUE" *) wire n7914_o;
  (* KEEP="TRUE" *) wire n7915_o;
  (* KEEP="TRUE" *) wire n7916_o;
  (* KEEP="TRUE" *) wire n7918_o;
  (* KEEP="TRUE" *) wire n7922_o;
  (* KEEP="TRUE" *) wire n7923_o;
  (* KEEP="TRUE" *) wire n7925_o;
  (* KEEP="TRUE" *) wire n7926_o;
  (* KEEP="TRUE" *) wire n7927_o;
  (* KEEP="TRUE" *) wire n7929_o;
  (* KEEP="TRUE" *) wire n7930_o;
  (* KEEP="TRUE" *) wire n7932_o;
  (* KEEP="TRUE" *) wire n7933_o;
  (* KEEP="TRUE" *) wire n7934_o;
  (* KEEP="TRUE" *) wire n7936_o;
  (* KEEP="TRUE" *) wire n7940_o;
  (* KEEP="TRUE" *) wire n7941_o;
  (* KEEP="TRUE" *) wire n7943_o;
  (* KEEP="TRUE" *) wire n7944_o;
  (* KEEP="TRUE" *) wire n7945_o;
  (* KEEP="TRUE" *) wire n7947_o;
  (* KEEP="TRUE" *) wire n7948_o;
  (* KEEP="TRUE" *) wire n7950_o;
  (* KEEP="TRUE" *) wire n7951_o;
  (* KEEP="TRUE" *) wire n7952_o;
  (* KEEP="TRUE" *) wire n7954_o;
  (* KEEP="TRUE" *) wire n7958_o;
  (* KEEP="TRUE" *) wire n7959_o;
  (* KEEP="TRUE" *) wire n7961_o;
  (* KEEP="TRUE" *) wire n7962_o;
  (* KEEP="TRUE" *) wire n7963_o;
  (* KEEP="TRUE" *) wire n7965_o;
  (* KEEP="TRUE" *) wire n7966_o;
  (* KEEP="TRUE" *) wire n7968_o;
  (* KEEP="TRUE" *) wire n7969_o;
  (* KEEP="TRUE" *) wire n7970_o;
  (* KEEP="TRUE" *) wire n7972_o;
  (* KEEP="TRUE" *) wire n7976_o;
  (* KEEP="TRUE" *) wire n7977_o;
  (* KEEP="TRUE" *) wire n7979_o;
  (* KEEP="TRUE" *) wire n7980_o;
  (* KEEP="TRUE" *) wire n7981_o;
  (* KEEP="TRUE" *) wire n7983_o;
  (* KEEP="TRUE" *) wire n7984_o;
  (* KEEP="TRUE" *) wire n7986_o;
  (* KEEP="TRUE" *) wire n7987_o;
  (* KEEP="TRUE" *) wire n7988_o;
  (* KEEP="TRUE" *) wire n7990_o;
  (* KEEP="TRUE" *) wire n7994_o;
  (* KEEP="TRUE" *) wire n7995_o;
  (* KEEP="TRUE" *) wire n7997_o;
  (* KEEP="TRUE" *) wire n7998_o;
  (* KEEP="TRUE" *) wire n7999_o;
  (* KEEP="TRUE" *) wire n8001_o;
  (* KEEP="TRUE" *) wire n8002_o;
  (* KEEP="TRUE" *) wire n8004_o;
  (* KEEP="TRUE" *) wire n8005_o;
  (* KEEP="TRUE" *) wire n8006_o;
  (* KEEP="TRUE" *) wire n8008_o;
  (* KEEP="TRUE" *) wire n8012_o;
  (* KEEP="TRUE" *) wire n8013_o;
  (* KEEP="TRUE" *) wire n8015_o;
  (* KEEP="TRUE" *) wire n8016_o;
  (* KEEP="TRUE" *) wire n8017_o;
  (* KEEP="TRUE" *) wire n8019_o;
  (* KEEP="TRUE" *) wire n8020_o;
  (* KEEP="TRUE" *) wire n8022_o;
  (* KEEP="TRUE" *) wire n8023_o;
  (* KEEP="TRUE" *) wire n8024_o;
  (* KEEP="TRUE" *) wire n8026_o;
  (* KEEP="TRUE" *) wire n8030_o;
  (* KEEP="TRUE" *) wire n8031_o;
  (* KEEP="TRUE" *) wire n8033_o;
  (* KEEP="TRUE" *) wire n8034_o;
  (* KEEP="TRUE" *) wire n8035_o;
  (* KEEP="TRUE" *) wire n8037_o;
  (* KEEP="TRUE" *) wire n8038_o;
  (* KEEP="TRUE" *) wire n8040_o;
  (* KEEP="TRUE" *) wire n8041_o;
  (* KEEP="TRUE" *) wire n8042_o;
  (* KEEP="TRUE" *) wire n8044_o;
  (* KEEP="TRUE" *) wire n8048_o;
  (* KEEP="TRUE" *) wire n8049_o;
  (* KEEP="TRUE" *) wire n8051_o;
  (* KEEP="TRUE" *) wire n8052_o;
  (* KEEP="TRUE" *) wire n8053_o;
  (* KEEP="TRUE" *) wire n8055_o;
  (* KEEP="TRUE" *) wire n8056_o;
  (* KEEP="TRUE" *) wire n8058_o;
  (* KEEP="TRUE" *) wire n8059_o;
  (* KEEP="TRUE" *) wire n8060_o;
  (* KEEP="TRUE" *) wire n8062_o;
  (* KEEP="TRUE" *) wire n8066_o;
  (* KEEP="TRUE" *) wire n8067_o;
  (* KEEP="TRUE" *) wire n8069_o;
  (* KEEP="TRUE" *) wire n8070_o;
  (* KEEP="TRUE" *) wire n8071_o;
  (* KEEP="TRUE" *) wire n8073_o;
  (* KEEP="TRUE" *) wire n8074_o;
  (* KEEP="TRUE" *) wire n8076_o;
  (* KEEP="TRUE" *) wire n8077_o;
  (* KEEP="TRUE" *) wire n8078_o;
  (* KEEP="TRUE" *) wire n8080_o;
  (* KEEP="TRUE" *) wire n8084_o;
  (* KEEP="TRUE" *) wire n8085_o;
  (* KEEP="TRUE" *) wire n8087_o;
  (* KEEP="TRUE" *) wire n8088_o;
  (* KEEP="TRUE" *) wire n8089_o;
  (* KEEP="TRUE" *) wire n8091_o;
  (* KEEP="TRUE" *) wire n8092_o;
  (* KEEP="TRUE" *) wire n8094_o;
  (* KEEP="TRUE" *) wire n8095_o;
  (* KEEP="TRUE" *) wire n8096_o;
  (* KEEP="TRUE" *) wire n8098_o;
  (* KEEP="TRUE" *) wire n8102_o;
  (* KEEP="TRUE" *) wire n8103_o;
  (* KEEP="TRUE" *) wire n8105_o;
  (* KEEP="TRUE" *) wire n8106_o;
  (* KEEP="TRUE" *) wire n8107_o;
  (* KEEP="TRUE" *) wire n8109_o;
  (* KEEP="TRUE" *) wire n8110_o;
  (* KEEP="TRUE" *) wire n8112_o;
  (* KEEP="TRUE" *) wire n8113_o;
  (* KEEP="TRUE" *) wire n8114_o;
  (* KEEP="TRUE" *) wire n8116_o;
  (* KEEP="TRUE" *) wire n8120_o;
  (* KEEP="TRUE" *) wire n8121_o;
  (* KEEP="TRUE" *) wire n8123_o;
  (* KEEP="TRUE" *) wire n8124_o;
  (* KEEP="TRUE" *) wire n8125_o;
  (* KEEP="TRUE" *) wire n8127_o;
  (* KEEP="TRUE" *) wire n8128_o;
  (* KEEP="TRUE" *) wire n8130_o;
  (* KEEP="TRUE" *) wire n8131_o;
  (* KEEP="TRUE" *) wire n8132_o;
  (* KEEP="TRUE" *) wire n8134_o;
  (* KEEP="TRUE" *) wire n8138_o;
  (* KEEP="TRUE" *) wire n8139_o;
  (* KEEP="TRUE" *) wire n8141_o;
  (* KEEP="TRUE" *) wire n8142_o;
  (* KEEP="TRUE" *) wire n8143_o;
  (* KEEP="TRUE" *) wire n8145_o;
  (* KEEP="TRUE" *) wire n8146_o;
  (* KEEP="TRUE" *) wire n8148_o;
  (* KEEP="TRUE" *) wire n8149_o;
  (* KEEP="TRUE" *) wire n8150_o;
  (* KEEP="TRUE" *) wire n8152_o;
  (* KEEP="TRUE" *) wire n8156_o;
  (* KEEP="TRUE" *) wire n8157_o;
  (* KEEP="TRUE" *) wire n8159_o;
  (* KEEP="TRUE" *) wire n8160_o;
  (* KEEP="TRUE" *) wire n8161_o;
  (* KEEP="TRUE" *) wire n8163_o;
  (* KEEP="TRUE" *) wire n8164_o;
  (* KEEP="TRUE" *) wire n8166_o;
  (* KEEP="TRUE" *) wire n8167_o;
  (* KEEP="TRUE" *) wire n8168_o;
  (* KEEP="TRUE" *) wire n8170_o;
  (* KEEP="TRUE" *) wire n8174_o;
  (* KEEP="TRUE" *) wire n8175_o;
  (* KEEP="TRUE" *) wire n8177_o;
  (* KEEP="TRUE" *) wire n8178_o;
  (* KEEP="TRUE" *) wire n8179_o;
  (* KEEP="TRUE" *) wire n8181_o;
  (* KEEP="TRUE" *) wire n8182_o;
  (* KEEP="TRUE" *) wire n8184_o;
  (* KEEP="TRUE" *) wire n8185_o;
  (* KEEP="TRUE" *) wire n8186_o;
  (* KEEP="TRUE" *) wire n8188_o;
  (* KEEP="TRUE" *) wire n8192_o;
  (* KEEP="TRUE" *) wire n8193_o;
  (* KEEP="TRUE" *) wire n8195_o;
  (* KEEP="TRUE" *) wire n8196_o;
  (* KEEP="TRUE" *) wire n8197_o;
  (* KEEP="TRUE" *) wire n8199_o;
  (* KEEP="TRUE" *) wire n8200_o;
  (* KEEP="TRUE" *) wire n8202_o;
  (* KEEP="TRUE" *) wire n8203_o;
  (* KEEP="TRUE" *) wire n8204_o;
  (* KEEP="TRUE" *) wire n8206_o;
  (* KEEP="TRUE" *) wire n8210_o;
  (* KEEP="TRUE" *) wire n8211_o;
  (* KEEP="TRUE" *) wire n8213_o;
  (* KEEP="TRUE" *) wire n8214_o;
  (* KEEP="TRUE" *) wire n8215_o;
  (* KEEP="TRUE" *) wire n8217_o;
  (* KEEP="TRUE" *) wire n8218_o;
  (* KEEP="TRUE" *) wire n8220_o;
  (* KEEP="TRUE" *) wire n8221_o;
  (* KEEP="TRUE" *) wire n8222_o;
  (* KEEP="TRUE" *) wire n8224_o;
  (* KEEP="TRUE" *) wire n8228_o;
  (* KEEP="TRUE" *) wire n8229_o;
  (* KEEP="TRUE" *) wire n8231_o;
  (* KEEP="TRUE" *) wire n8232_o;
  (* KEEP="TRUE" *) wire n8233_o;
  (* KEEP="TRUE" *) wire n8235_o;
  (* KEEP="TRUE" *) wire n8236_o;
  (* KEEP="TRUE" *) wire n8238_o;
  (* KEEP="TRUE" *) wire n8239_o;
  (* KEEP="TRUE" *) wire n8240_o;
  (* KEEP="TRUE" *) wire n8242_o;
  (* KEEP="TRUE" *) wire n8246_o;
  (* KEEP="TRUE" *) wire n8247_o;
  (* KEEP="TRUE" *) wire n8249_o;
  (* KEEP="TRUE" *) wire n8250_o;
  (* KEEP="TRUE" *) wire n8251_o;
  (* KEEP="TRUE" *) wire n8253_o;
  (* KEEP="TRUE" *) wire n8254_o;
  (* KEEP="TRUE" *) wire n8256_o;
  (* KEEP="TRUE" *) wire n8257_o;
  (* KEEP="TRUE" *) wire n8258_o;
  (* KEEP="TRUE" *) wire n8260_o;
  (* KEEP="TRUE" *) wire n8264_o;
  (* KEEP="TRUE" *) wire n8265_o;
  (* KEEP="TRUE" *) wire n8267_o;
  (* KEEP="TRUE" *) wire n8268_o;
  (* KEEP="TRUE" *) wire n8269_o;
  (* KEEP="TRUE" *) wire n8271_o;
  (* KEEP="TRUE" *) wire n8272_o;
  (* KEEP="TRUE" *) wire n8274_o;
  (* KEEP="TRUE" *) wire n8275_o;
  (* KEEP="TRUE" *) wire n8276_o;
  (* KEEP="TRUE" *) wire n8278_o;
  (* KEEP="TRUE" *) wire n8282_o;
  (* KEEP="TRUE" *) wire n8283_o;
  (* KEEP="TRUE" *) wire n8285_o;
  (* KEEP="TRUE" *) wire n8286_o;
  (* KEEP="TRUE" *) wire n8287_o;
  (* KEEP="TRUE" *) wire n8289_o;
  (* KEEP="TRUE" *) wire n8290_o;
  (* KEEP="TRUE" *) wire n8292_o;
  (* KEEP="TRUE" *) wire n8293_o;
  (* KEEP="TRUE" *) wire n8294_o;
  (* KEEP="TRUE" *) wire n8296_o;
  (* KEEP="TRUE" *) wire n8300_o;
  (* KEEP="TRUE" *) wire n8301_o;
  (* KEEP="TRUE" *) wire n8303_o;
  (* KEEP="TRUE" *) wire n8304_o;
  (* KEEP="TRUE" *) wire n8305_o;
  (* KEEP="TRUE" *) wire n8307_o;
  (* KEEP="TRUE" *) wire n8308_o;
  (* KEEP="TRUE" *) wire n8310_o;
  (* KEEP="TRUE" *) wire n8311_o;
  (* KEEP="TRUE" *) wire n8312_o;
  (* KEEP="TRUE" *) wire n8314_o;
  (* KEEP="TRUE" *) wire n8318_o;
  (* KEEP="TRUE" *) wire n8319_o;
  (* KEEP="TRUE" *) wire n8321_o;
  (* KEEP="TRUE" *) wire n8322_o;
  (* KEEP="TRUE" *) wire n8323_o;
  (* KEEP="TRUE" *) wire n8325_o;
  (* KEEP="TRUE" *) wire n8326_o;
  (* KEEP="TRUE" *) wire n8328_o;
  (* KEEP="TRUE" *) wire n8329_o;
  (* KEEP="TRUE" *) wire n8330_o;
  (* KEEP="TRUE" *) wire n8332_o;
  (* KEEP="TRUE" *) wire n8336_o;
  (* KEEP="TRUE" *) wire n8337_o;
  (* KEEP="TRUE" *) wire n8339_o;
  (* KEEP="TRUE" *) wire n8340_o;
  (* KEEP="TRUE" *) wire n8341_o;
  (* KEEP="TRUE" *) wire n8343_o;
  (* KEEP="TRUE" *) wire n8344_o;
  (* KEEP="TRUE" *) wire n8346_o;
  (* KEEP="TRUE" *) wire n8347_o;
  (* KEEP="TRUE" *) wire n8348_o;
  (* KEEP="TRUE" *) wire n8350_o;
  (* KEEP="TRUE" *) wire n8354_o;
  (* KEEP="TRUE" *) wire n8355_o;
  (* KEEP="TRUE" *) wire n8357_o;
  (* KEEP="TRUE" *) wire n8358_o;
  (* KEEP="TRUE" *) wire n8359_o;
  (* KEEP="TRUE" *) wire n8361_o;
  (* KEEP="TRUE" *) wire n8362_o;
  (* KEEP="TRUE" *) wire n8364_o;
  (* KEEP="TRUE" *) wire n8365_o;
  (* KEEP="TRUE" *) wire n8366_o;
  (* KEEP="TRUE" *) wire n8368_o;
  (* KEEP="TRUE" *) wire n8372_o;
  (* KEEP="TRUE" *) wire n8373_o;
  (* KEEP="TRUE" *) wire n8375_o;
  (* KEEP="TRUE" *) wire n8376_o;
  (* KEEP="TRUE" *) wire n8377_o;
  (* KEEP="TRUE" *) wire n8379_o;
  (* KEEP="TRUE" *) wire n8380_o;
  (* KEEP="TRUE" *) wire n8382_o;
  (* KEEP="TRUE" *) wire n8383_o;
  (* KEEP="TRUE" *) wire n8384_o;
  (* KEEP="TRUE" *) wire n8386_o;
  (* KEEP="TRUE" *) wire n8390_o;
  (* KEEP="TRUE" *) wire n8391_o;
  (* KEEP="TRUE" *) wire n8393_o;
  (* KEEP="TRUE" *) wire n8394_o;
  (* KEEP="TRUE" *) wire n8395_o;
  (* KEEP="TRUE" *) wire n8397_o;
  (* KEEP="TRUE" *) wire n8398_o;
  (* KEEP="TRUE" *) wire n8400_o;
  (* KEEP="TRUE" *) wire n8401_o;
  (* KEEP="TRUE" *) wire n8402_o;
  (* KEEP="TRUE" *) wire n8404_o;
  (* KEEP="TRUE" *) wire n8408_o;
  (* KEEP="TRUE" *) wire n8409_o;
  (* KEEP="TRUE" *) wire n8411_o;
  (* KEEP="TRUE" *) wire n8412_o;
  (* KEEP="TRUE" *) wire n8413_o;
  (* KEEP="TRUE" *) wire n8415_o;
  (* KEEP="TRUE" *) wire n8416_o;
  (* KEEP="TRUE" *) wire n8418_o;
  (* KEEP="TRUE" *) wire n8419_o;
  (* KEEP="TRUE" *) wire n8420_o;
  (* KEEP="TRUE" *) wire n8422_o;
  (* KEEP="TRUE" *) wire n8426_o;
  (* KEEP="TRUE" *) wire n8427_o;
  (* KEEP="TRUE" *) wire n8429_o;
  (* KEEP="TRUE" *) wire n8430_o;
  (* KEEP="TRUE" *) wire n8431_o;
  (* KEEP="TRUE" *) wire n8433_o;
  (* KEEP="TRUE" *) wire n8434_o;
  (* KEEP="TRUE" *) wire n8436_o;
  (* KEEP="TRUE" *) wire n8437_o;
  (* KEEP="TRUE" *) wire n8438_o;
  (* KEEP="TRUE" *) wire n8440_o;
  (* KEEP="TRUE" *) wire n8444_o;
  (* KEEP="TRUE" *) wire n8445_o;
  (* KEEP="TRUE" *) wire n8447_o;
  (* KEEP="TRUE" *) wire n8448_o;
  (* KEEP="TRUE" *) wire n8449_o;
  (* KEEP="TRUE" *) wire n8451_o;
  (* KEEP="TRUE" *) wire n8452_o;
  (* KEEP="TRUE" *) wire n8454_o;
  (* KEEP="TRUE" *) wire n8455_o;
  (* KEEP="TRUE" *) wire n8456_o;
  (* KEEP="TRUE" *) wire n8458_o;
  (* KEEP="TRUE" *) wire n8462_o;
  (* KEEP="TRUE" *) wire n8463_o;
  (* KEEP="TRUE" *) wire n8465_o;
  (* KEEP="TRUE" *) wire n8466_o;
  (* KEEP="TRUE" *) wire n8467_o;
  (* KEEP="TRUE" *) wire n8469_o;
  (* KEEP="TRUE" *) wire n8470_o;
  (* KEEP="TRUE" *) wire n8472_o;
  (* KEEP="TRUE" *) wire n8473_o;
  (* KEEP="TRUE" *) wire n8474_o;
  (* KEEP="TRUE" *) wire n8476_o;
  (* KEEP="TRUE" *) wire n8480_o;
  (* KEEP="TRUE" *) wire n8481_o;
  (* KEEP="TRUE" *) wire n8483_o;
  (* KEEP="TRUE" *) wire n8484_o;
  (* KEEP="TRUE" *) wire n8485_o;
  (* KEEP="TRUE" *) wire n8487_o;
  (* KEEP="TRUE" *) wire n8488_o;
  (* KEEP="TRUE" *) wire n8490_o;
  (* KEEP="TRUE" *) wire n8491_o;
  (* KEEP="TRUE" *) wire n8492_o;
  (* KEEP="TRUE" *) wire n8494_o;
  (* KEEP="TRUE" *) wire n8498_o;
  (* KEEP="TRUE" *) wire n8499_o;
  (* KEEP="TRUE" *) wire n8501_o;
  (* KEEP="TRUE" *) wire n8502_o;
  (* KEEP="TRUE" *) wire n8503_o;
  (* KEEP="TRUE" *) wire n8505_o;
  (* KEEP="TRUE" *) wire n8506_o;
  (* KEEP="TRUE" *) wire n8508_o;
  (* KEEP="TRUE" *) wire n8509_o;
  (* KEEP="TRUE" *) wire n8510_o;
  (* KEEP="TRUE" *) wire n8512_o;
  (* KEEP="TRUE" *) wire n8516_o;
  (* KEEP="TRUE" *) wire n8517_o;
  (* KEEP="TRUE" *) wire n8519_o;
  (* KEEP="TRUE" *) wire n8520_o;
  (* KEEP="TRUE" *) wire n8521_o;
  (* KEEP="TRUE" *) wire n8523_o;
  (* KEEP="TRUE" *) wire n8524_o;
  (* KEEP="TRUE" *) wire n8526_o;
  (* KEEP="TRUE" *) wire n8527_o;
  (* KEEP="TRUE" *) wire n8528_o;
  (* KEEP="TRUE" *) wire n8530_o;
  (* KEEP="TRUE" *) wire n8534_o;
  (* KEEP="TRUE" *) wire n8535_o;
  (* KEEP="TRUE" *) wire n8537_o;
  (* KEEP="TRUE" *) wire n8538_o;
  (* KEEP="TRUE" *) wire n8539_o;
  (* KEEP="TRUE" *) wire n8541_o;
  (* KEEP="TRUE" *) wire n8542_o;
  (* KEEP="TRUE" *) wire n8544_o;
  (* KEEP="TRUE" *) wire n8545_o;
  (* KEEP="TRUE" *) wire n8546_o;
  (* KEEP="TRUE" *) wire n8548_o;
  (* KEEP="TRUE" *) wire n8552_o;
  (* KEEP="TRUE" *) wire n8553_o;
  (* KEEP="TRUE" *) wire n8555_o;
  (* KEEP="TRUE" *) wire n8556_o;
  (* KEEP="TRUE" *) wire n8557_o;
  (* KEEP="TRUE" *) wire n8559_o;
  (* KEEP="TRUE" *) wire n8560_o;
  (* KEEP="TRUE" *) wire n8562_o;
  (* KEEP="TRUE" *) wire n8563_o;
  (* KEEP="TRUE" *) wire n8564_o;
  (* KEEP="TRUE" *) wire n8566_o;
  (* KEEP="TRUE" *) wire n8570_o;
  (* KEEP="TRUE" *) wire n8571_o;
  (* KEEP="TRUE" *) wire n8573_o;
  (* KEEP="TRUE" *) wire n8574_o;
  (* KEEP="TRUE" *) wire n8575_o;
  (* KEEP="TRUE" *) wire n8577_o;
  (* KEEP="TRUE" *) wire n8578_o;
  (* KEEP="TRUE" *) wire n8580_o;
  (* KEEP="TRUE" *) wire n8581_o;
  (* KEEP="TRUE" *) wire n8582_o;
  (* KEEP="TRUE" *) wire n8584_o;
  (* KEEP="TRUE" *) wire n8588_o;
  (* KEEP="TRUE" *) wire n8589_o;
  (* KEEP="TRUE" *) wire n8591_o;
  (* KEEP="TRUE" *) wire n8592_o;
  (* KEEP="TRUE" *) wire n8593_o;
  (* KEEP="TRUE" *) wire n8595_o;
  (* KEEP="TRUE" *) wire n8596_o;
  (* KEEP="TRUE" *) wire n8598_o;
  (* KEEP="TRUE" *) wire n8599_o;
  (* KEEP="TRUE" *) wire n8600_o;
  (* KEEP="TRUE" *) wire n8602_o;
  (* KEEP="TRUE" *) wire n8606_o;
  (* KEEP="TRUE" *) wire n8607_o;
  (* KEEP="TRUE" *) wire n8609_o;
  (* KEEP="TRUE" *) wire n8610_o;
  (* KEEP="TRUE" *) wire n8611_o;
  (* KEEP="TRUE" *) wire n8613_o;
  (* KEEP="TRUE" *) wire n8614_o;
  (* KEEP="TRUE" *) wire n8616_o;
  (* KEEP="TRUE" *) wire n8617_o;
  (* KEEP="TRUE" *) wire n8618_o;
  (* KEEP="TRUE" *) wire n8620_o;
  (* KEEP="TRUE" *) wire n8624_o;
  (* KEEP="TRUE" *) wire n8625_o;
  (* KEEP="TRUE" *) wire n8627_o;
  (* KEEP="TRUE" *) wire n8628_o;
  (* KEEP="TRUE" *) wire n8629_o;
  (* KEEP="TRUE" *) wire n8631_o;
  (* KEEP="TRUE" *) wire n8632_o;
  (* KEEP="TRUE" *) wire n8634_o;
  (* KEEP="TRUE" *) wire n8635_o;
  (* KEEP="TRUE" *) wire n8636_o;
  (* KEEP="TRUE" *) wire n8638_o;
  (* KEEP="TRUE" *) wire n8642_o;
  (* KEEP="TRUE" *) wire n8643_o;
  (* KEEP="TRUE" *) wire n8645_o;
  (* KEEP="TRUE" *) wire n8646_o;
  (* KEEP="TRUE" *) wire n8647_o;
  (* KEEP="TRUE" *) wire n8649_o;
  (* KEEP="TRUE" *) wire n8650_o;
  (* KEEP="TRUE" *) wire n8652_o;
  (* KEEP="TRUE" *) wire n8653_o;
  (* KEEP="TRUE" *) wire n8654_o;
  (* KEEP="TRUE" *) wire n8656_o;
  (* KEEP="TRUE" *) wire n8660_o;
  (* KEEP="TRUE" *) wire n8661_o;
  (* KEEP="TRUE" *) wire n8663_o;
  (* KEEP="TRUE" *) wire n8664_o;
  (* KEEP="TRUE" *) wire n8665_o;
  (* KEEP="TRUE" *) wire n8667_o;
  (* KEEP="TRUE" *) wire n8668_o;
  (* KEEP="TRUE" *) wire n8670_o;
  (* KEEP="TRUE" *) wire n8671_o;
  (* KEEP="TRUE" *) wire n8672_o;
  (* KEEP="TRUE" *) wire n8674_o;
  (* KEEP="TRUE" *) wire n8678_o;
  (* KEEP="TRUE" *) wire n8679_o;
  (* KEEP="TRUE" *) wire n8681_o;
  (* KEEP="TRUE" *) wire n8682_o;
  (* KEEP="TRUE" *) wire n8683_o;
  (* KEEP="TRUE" *) wire n8685_o;
  (* KEEP="TRUE" *) wire n8686_o;
  (* KEEP="TRUE" *) wire n8688_o;
  (* KEEP="TRUE" *) wire n8689_o;
  (* KEEP="TRUE" *) wire n8690_o;
  (* KEEP="TRUE" *) wire n8692_o;
  (* KEEP="TRUE" *) wire n8696_o;
  (* KEEP="TRUE" *) wire n8697_o;
  (* KEEP="TRUE" *) wire n8699_o;
  (* KEEP="TRUE" *) wire n8700_o;
  (* KEEP="TRUE" *) wire n8701_o;
  (* KEEP="TRUE" *) wire n8703_o;
  (* KEEP="TRUE" *) wire n8704_o;
  (* KEEP="TRUE" *) wire n8706_o;
  (* KEEP="TRUE" *) wire n8707_o;
  (* KEEP="TRUE" *) wire n8708_o;
  (* KEEP="TRUE" *) wire n8710_o;
  (* KEEP="TRUE" *) wire n8714_o;
  (* KEEP="TRUE" *) wire n8715_o;
  (* KEEP="TRUE" *) wire n8717_o;
  (* KEEP="TRUE" *) wire n8718_o;
  (* KEEP="TRUE" *) wire n8719_o;
  (* KEEP="TRUE" *) wire n8721_o;
  (* KEEP="TRUE" *) wire n8722_o;
  (* KEEP="TRUE" *) wire n8724_o;
  (* KEEP="TRUE" *) wire n8725_o;
  (* KEEP="TRUE" *) wire n8726_o;
  (* KEEP="TRUE" *) wire n8728_o;
  (* KEEP="TRUE" *) wire n8732_o;
  (* KEEP="TRUE" *) wire n8733_o;
  (* KEEP="TRUE" *) wire n8735_o;
  (* KEEP="TRUE" *) wire n8736_o;
  (* KEEP="TRUE" *) wire n8737_o;
  (* KEEP="TRUE" *) wire n8739_o;
  (* KEEP="TRUE" *) wire n8740_o;
  (* KEEP="TRUE" *) wire n8742_o;
  (* KEEP="TRUE" *) wire n8743_o;
  (* KEEP="TRUE" *) wire n8744_o;
  (* KEEP="TRUE" *) wire n8746_o;
  (* KEEP="TRUE" *) wire n8750_o;
  (* KEEP="TRUE" *) wire n8751_o;
  (* KEEP="TRUE" *) wire n8753_o;
  (* KEEP="TRUE" *) wire n8754_o;
  (* KEEP="TRUE" *) wire n8755_o;
  (* KEEP="TRUE" *) wire n8757_o;
  (* KEEP="TRUE" *) wire n8758_o;
  (* KEEP="TRUE" *) wire n8760_o;
  (* KEEP="TRUE" *) wire n8761_o;
  (* KEEP="TRUE" *) wire n8762_o;
  (* KEEP="TRUE" *) wire n8764_o;
  (* KEEP="TRUE" *) wire n8768_o;
  (* KEEP="TRUE" *) wire n8769_o;
  (* KEEP="TRUE" *) wire n8771_o;
  (* KEEP="TRUE" *) wire n8772_o;
  (* KEEP="TRUE" *) wire n8773_o;
  (* KEEP="TRUE" *) wire n8775_o;
  (* KEEP="TRUE" *) wire n8776_o;
  (* KEEP="TRUE" *) wire n8778_o;
  (* KEEP="TRUE" *) wire n8779_o;
  (* KEEP="TRUE" *) wire n8780_o;
  (* KEEP="TRUE" *) wire n8782_o;
  (* KEEP="TRUE" *) wire n8786_o;
  (* KEEP="TRUE" *) wire n8787_o;
  (* KEEP="TRUE" *) wire n8789_o;
  (* KEEP="TRUE" *) wire n8790_o;
  (* KEEP="TRUE" *) wire n8791_o;
  (* KEEP="TRUE" *) wire n8793_o;
  (* KEEP="TRUE" *) wire n8794_o;
  (* KEEP="TRUE" *) wire n8796_o;
  (* KEEP="TRUE" *) wire n8797_o;
  (* KEEP="TRUE" *) wire n8798_o;
  (* KEEP="TRUE" *) wire n8800_o;
  (* KEEP="TRUE" *) wire n8804_o;
  (* KEEP="TRUE" *) wire n8805_o;
  (* KEEP="TRUE" *) wire n8807_o;
  (* KEEP="TRUE" *) wire n8808_o;
  (* KEEP="TRUE" *) wire n8809_o;
  (* KEEP="TRUE" *) wire n8811_o;
  (* KEEP="TRUE" *) wire n8812_o;
  (* KEEP="TRUE" *) wire n8814_o;
  (* KEEP="TRUE" *) wire n8815_o;
  (* KEEP="TRUE" *) wire n8816_o;
  (* KEEP="TRUE" *) wire n8818_o;
  (* KEEP="TRUE" *) wire n8822_o;
  (* KEEP="TRUE" *) wire n8823_o;
  (* KEEP="TRUE" *) wire n8825_o;
  (* KEEP="TRUE" *) wire n8826_o;
  (* KEEP="TRUE" *) wire n8827_o;
  (* KEEP="TRUE" *) wire n8829_o;
  (* KEEP="TRUE" *) wire n8830_o;
  (* KEEP="TRUE" *) wire n8832_o;
  (* KEEP="TRUE" *) wire n8833_o;
  (* KEEP="TRUE" *) wire n8834_o;
  (* KEEP="TRUE" *) wire n8836_o;
  (* KEEP="TRUE" *) wire n8840_o;
  (* KEEP="TRUE" *) wire n8841_o;
  (* KEEP="TRUE" *) wire n8843_o;
  (* KEEP="TRUE" *) wire n8844_o;
  (* KEEP="TRUE" *) wire n8845_o;
  (* KEEP="TRUE" *) wire n8847_o;
  (* KEEP="TRUE" *) wire n8848_o;
  (* KEEP="TRUE" *) wire n8850_o;
  (* KEEP="TRUE" *) wire n8851_o;
  (* KEEP="TRUE" *) wire n8852_o;
  (* KEEP="TRUE" *) wire n8854_o;
  (* KEEP="TRUE" *) wire n8858_o;
  (* KEEP="TRUE" *) wire n8859_o;
  (* KEEP="TRUE" *) wire n8861_o;
  (* KEEP="TRUE" *) wire n8862_o;
  (* KEEP="TRUE" *) wire n8863_o;
  (* KEEP="TRUE" *) wire n8865_o;
  (* KEEP="TRUE" *) wire n8866_o;
  (* KEEP="TRUE" *) wire n8868_o;
  (* KEEP="TRUE" *) wire n8869_o;
  (* KEEP="TRUE" *) wire n8870_o;
  (* KEEP="TRUE" *) wire n8872_o;
  (* KEEP="TRUE" *) wire n8876_o;
  (* KEEP="TRUE" *) wire n8877_o;
  (* KEEP="TRUE" *) wire n8879_o;
  (* KEEP="TRUE" *) wire n8880_o;
  (* KEEP="TRUE" *) wire n8881_o;
  (* KEEP="TRUE" *) wire n8883_o;
  (* KEEP="TRUE" *) wire n8884_o;
  (* KEEP="TRUE" *) wire n8886_o;
  (* KEEP="TRUE" *) wire n8887_o;
  (* KEEP="TRUE" *) wire n8888_o;
  (* KEEP="TRUE" *) wire n8890_o;
  (* KEEP="TRUE" *) wire n8894_o;
  (* KEEP="TRUE" *) wire n8895_o;
  (* KEEP="TRUE" *) wire n8897_o;
  (* KEEP="TRUE" *) wire n8898_o;
  (* KEEP="TRUE" *) wire n8899_o;
  (* KEEP="TRUE" *) wire n8901_o;
  (* KEEP="TRUE" *) wire n8902_o;
  (* KEEP="TRUE" *) wire n8904_o;
  (* KEEP="TRUE" *) wire n8905_o;
  (* KEEP="TRUE" *) wire n8906_o;
  (* KEEP="TRUE" *) wire n8908_o;
  (* KEEP="TRUE" *) wire n8912_o;
  (* KEEP="TRUE" *) wire n8913_o;
  (* KEEP="TRUE" *) wire n8915_o;
  (* KEEP="TRUE" *) wire n8916_o;
  (* KEEP="TRUE" *) wire n8917_o;
  (* KEEP="TRUE" *) wire n8919_o;
  (* KEEP="TRUE" *) wire n8920_o;
  (* KEEP="TRUE" *) wire n8922_o;
  (* KEEP="TRUE" *) wire n8923_o;
  (* KEEP="TRUE" *) wire n8924_o;
  (* KEEP="TRUE" *) wire n8926_o;
  (* KEEP="TRUE" *) wire n8930_o;
  (* KEEP="TRUE" *) wire n8931_o;
  (* KEEP="TRUE" *) wire n8933_o;
  (* KEEP="TRUE" *) wire n8934_o;
  (* KEEP="TRUE" *) wire n8935_o;
  (* KEEP="TRUE" *) wire n8937_o;
  (* KEEP="TRUE" *) wire n8938_o;
  (* KEEP="TRUE" *) wire n8940_o;
  (* KEEP="TRUE" *) wire n8941_o;
  (* KEEP="TRUE" *) wire n8942_o;
  (* KEEP="TRUE" *) wire n8944_o;
  (* KEEP="TRUE" *) wire n8948_o;
  (* KEEP="TRUE" *) wire n8949_o;
  (* KEEP="TRUE" *) wire n8951_o;
  (* KEEP="TRUE" *) wire n8952_o;
  (* KEEP="TRUE" *) wire n8953_o;
  (* KEEP="TRUE" *) wire n8955_o;
  (* KEEP="TRUE" *) wire n8956_o;
  (* KEEP="TRUE" *) wire n8958_o;
  (* KEEP="TRUE" *) wire n8959_o;
  (* KEEP="TRUE" *) wire n8960_o;
  (* KEEP="TRUE" *) wire n8962_o;
  (* KEEP="TRUE" *) wire n8966_o;
  (* KEEP="TRUE" *) wire n8967_o;
  (* KEEP="TRUE" *) wire n8969_o;
  (* KEEP="TRUE" *) wire n8970_o;
  (* KEEP="TRUE" *) wire n8971_o;
  (* KEEP="TRUE" *) wire n8973_o;
  (* KEEP="TRUE" *) wire n8974_o;
  (* KEEP="TRUE" *) wire n8976_o;
  (* KEEP="TRUE" *) wire n8977_o;
  (* KEEP="TRUE" *) wire n8978_o;
  (* KEEP="TRUE" *) wire n8980_o;
  (* KEEP="TRUE" *) wire n8984_o;
  (* KEEP="TRUE" *) wire n8985_o;
  (* KEEP="TRUE" *) wire n8987_o;
  (* KEEP="TRUE" *) wire n8988_o;
  (* KEEP="TRUE" *) wire n8989_o;
  (* KEEP="TRUE" *) wire n8991_o;
  (* KEEP="TRUE" *) wire n8992_o;
  (* KEEP="TRUE" *) wire n8994_o;
  (* KEEP="TRUE" *) wire n8995_o;
  (* KEEP="TRUE" *) wire n8996_o;
  (* KEEP="TRUE" *) wire n8998_o;
  (* KEEP="TRUE" *) wire n9002_o;
  (* KEEP="TRUE" *) wire n9003_o;
  (* KEEP="TRUE" *) wire n9005_o;
  (* KEEP="TRUE" *) wire n9006_o;
  (* KEEP="TRUE" *) wire n9007_o;
  (* KEEP="TRUE" *) wire n9009_o;
  (* KEEP="TRUE" *) wire n9010_o;
  (* KEEP="TRUE" *) wire n9012_o;
  (* KEEP="TRUE" *) wire n9013_o;
  (* KEEP="TRUE" *) wire n9014_o;
  (* KEEP="TRUE" *) wire n9016_o;
  (* KEEP="TRUE" *) wire n9020_o;
  (* KEEP="TRUE" *) wire n9021_o;
  (* KEEP="TRUE" *) wire n9023_o;
  (* KEEP="TRUE" *) wire n9024_o;
  (* KEEP="TRUE" *) wire n9025_o;
  (* KEEP="TRUE" *) wire n9027_o;
  (* KEEP="TRUE" *) wire n9028_o;
  (* KEEP="TRUE" *) wire n9030_o;
  (* KEEP="TRUE" *) wire n9031_o;
  (* KEEP="TRUE" *) wire n9032_o;
  (* KEEP="TRUE" *) wire n9034_o;
  (* KEEP="TRUE" *) wire n9038_o;
  (* KEEP="TRUE" *) wire n9039_o;
  (* KEEP="TRUE" *) wire n9041_o;
  (* KEEP="TRUE" *) wire n9042_o;
  (* KEEP="TRUE" *) wire n9043_o;
  (* KEEP="TRUE" *) wire n9045_o;
  (* KEEP="TRUE" *) wire n9046_o;
  (* KEEP="TRUE" *) wire n9048_o;
  (* KEEP="TRUE" *) wire n9049_o;
  (* KEEP="TRUE" *) wire n9050_o;
  (* KEEP="TRUE" *) wire n9052_o;
  (* KEEP="TRUE" *) wire n9056_o;
  (* KEEP="TRUE" *) wire n9057_o;
  (* KEEP="TRUE" *) wire n9059_o;
  (* KEEP="TRUE" *) wire n9060_o;
  (* KEEP="TRUE" *) wire n9061_o;
  (* KEEP="TRUE" *) wire n9063_o;
  (* KEEP="TRUE" *) wire n9064_o;
  (* KEEP="TRUE" *) wire n9066_o;
  (* KEEP="TRUE" *) wire n9067_o;
  (* KEEP="TRUE" *) wire n9068_o;
  (* KEEP="TRUE" *) wire n9070_o;
  (* KEEP="TRUE" *) wire n9074_o;
  (* KEEP="TRUE" *) wire n9075_o;
  (* KEEP="TRUE" *) wire n9077_o;
  (* KEEP="TRUE" *) wire n9078_o;
  (* KEEP="TRUE" *) wire n9079_o;
  (* KEEP="TRUE" *) wire n9081_o;
  (* KEEP="TRUE" *) wire n9082_o;
  (* KEEP="TRUE" *) wire n9084_o;
  (* KEEP="TRUE" *) wire n9085_o;
  (* KEEP="TRUE" *) wire n9086_o;
  (* KEEP="TRUE" *) wire n9088_o;
  (* KEEP="TRUE" *) wire n9092_o;
  (* KEEP="TRUE" *) wire n9093_o;
  (* KEEP="TRUE" *) wire n9095_o;
  (* KEEP="TRUE" *) wire n9096_o;
  (* KEEP="TRUE" *) wire n9097_o;
  (* KEEP="TRUE" *) wire n9099_o;
  (* KEEP="TRUE" *) wire n9100_o;
  (* KEEP="TRUE" *) wire n9102_o;
  (* KEEP="TRUE" *) wire n9103_o;
  (* KEEP="TRUE" *) wire n9104_o;
  (* KEEP="TRUE" *) wire n9106_o;
  (* KEEP="TRUE" *) wire n9110_o;
  (* KEEP="TRUE" *) wire n9111_o;
  (* KEEP="TRUE" *) wire n9113_o;
  (* KEEP="TRUE" *) wire n9114_o;
  (* KEEP="TRUE" *) wire n9115_o;
  (* KEEP="TRUE" *) wire n9117_o;
  (* KEEP="TRUE" *) wire n9118_o;
  (* KEEP="TRUE" *) wire n9120_o;
  (* KEEP="TRUE" *) wire n9121_o;
  (* KEEP="TRUE" *) wire n9122_o;
  (* KEEP="TRUE" *) wire n9124_o;
  (* KEEP="TRUE" *) wire n9128_o;
  (* KEEP="TRUE" *) wire n9129_o;
  (* KEEP="TRUE" *) wire n9131_o;
  (* KEEP="TRUE" *) wire n9132_o;
  (* KEEP="TRUE" *) wire n9133_o;
  (* KEEP="TRUE" *) wire n9135_o;
  (* KEEP="TRUE" *) wire n9136_o;
  (* KEEP="TRUE" *) wire n9138_o;
  (* KEEP="TRUE" *) wire n9139_o;
  (* KEEP="TRUE" *) wire n9140_o;
  (* KEEP="TRUE" *) wire n9142_o;
  (* KEEP="TRUE" *) wire n9146_o;
  (* KEEP="TRUE" *) wire n9147_o;
  (* KEEP="TRUE" *) wire n9149_o;
  (* KEEP="TRUE" *) wire n9150_o;
  (* KEEP="TRUE" *) wire n9151_o;
  (* KEEP="TRUE" *) wire n9153_o;
  (* KEEP="TRUE" *) wire n9154_o;
  (* KEEP="TRUE" *) wire n9156_o;
  (* KEEP="TRUE" *) wire n9157_o;
  (* KEEP="TRUE" *) wire n9158_o;
  (* KEEP="TRUE" *) wire n9160_o;
  (* KEEP="TRUE" *) wire n9164_o;
  (* KEEP="TRUE" *) wire n9165_o;
  (* KEEP="TRUE" *) wire n9167_o;
  (* KEEP="TRUE" *) wire n9168_o;
  (* KEEP="TRUE" *) wire n9169_o;
  (* KEEP="TRUE" *) wire n9171_o;
  (* KEEP="TRUE" *) wire n9172_o;
  (* KEEP="TRUE" *) wire n9174_o;
  (* KEEP="TRUE" *) wire n9175_o;
  (* KEEP="TRUE" *) wire n9176_o;
  (* KEEP="TRUE" *) wire n9178_o;
  (* KEEP="TRUE" *) wire n9182_o;
  (* KEEP="TRUE" *) wire n9183_o;
  (* KEEP="TRUE" *) wire n9185_o;
  (* KEEP="TRUE" *) wire n9186_o;
  (* KEEP="TRUE" *) wire n9187_o;
  (* KEEP="TRUE" *) wire n9189_o;
  (* KEEP="TRUE" *) wire n9190_o;
  (* KEEP="TRUE" *) wire n9192_o;
  (* KEEP="TRUE" *) wire n9193_o;
  (* KEEP="TRUE" *) wire n9194_o;
  (* KEEP="TRUE" *) wire n9196_o;
  (* KEEP="TRUE" *) wire n9200_o;
  (* KEEP="TRUE" *) wire n9201_o;
  (* KEEP="TRUE" *) wire n9203_o;
  (* KEEP="TRUE" *) wire n9204_o;
  (* KEEP="TRUE" *) wire n9205_o;
  (* KEEP="TRUE" *) wire n9207_o;
  (* KEEP="TRUE" *) wire n9208_o;
  (* KEEP="TRUE" *) wire n9210_o;
  (* KEEP="TRUE" *) wire n9211_o;
  (* KEEP="TRUE" *) wire n9212_o;
  (* KEEP="TRUE" *) wire n9214_o;
  (* KEEP="TRUE" *) wire n9218_o;
  (* KEEP="TRUE" *) wire n9219_o;
  (* KEEP="TRUE" *) wire n9221_o;
  (* KEEP="TRUE" *) wire n9222_o;
  (* KEEP="TRUE" *) wire n9223_o;
  (* KEEP="TRUE" *) wire n9225_o;
  (* KEEP="TRUE" *) wire n9226_o;
  (* KEEP="TRUE" *) wire n9228_o;
  (* KEEP="TRUE" *) wire n9229_o;
  (* KEEP="TRUE" *) wire n9230_o;
  (* KEEP="TRUE" *) wire n9232_o;
  (* KEEP="TRUE" *) wire n9236_o;
  (* KEEP="TRUE" *) wire n9237_o;
  (* KEEP="TRUE" *) wire n9239_o;
  (* KEEP="TRUE" *) wire n9240_o;
  (* KEEP="TRUE" *) wire n9241_o;
  (* KEEP="TRUE" *) wire n9243_o;
  (* KEEP="TRUE" *) wire n9244_o;
  (* KEEP="TRUE" *) wire n9246_o;
  (* KEEP="TRUE" *) wire n9247_o;
  (* KEEP="TRUE" *) wire n9248_o;
  (* KEEP="TRUE" *) wire n9250_o;
  (* KEEP="TRUE" *) wire n9254_o;
  (* KEEP="TRUE" *) wire n9255_o;
  (* KEEP="TRUE" *) wire n9257_o;
  (* KEEP="TRUE" *) wire n9258_o;
  (* KEEP="TRUE" *) wire n9259_o;
  (* KEEP="TRUE" *) wire n9261_o;
  (* KEEP="TRUE" *) wire n9262_o;
  (* KEEP="TRUE" *) wire n9264_o;
  (* KEEP="TRUE" *) wire n9265_o;
  (* KEEP="TRUE" *) wire n9266_o;
  (* KEEP="TRUE" *) wire n9268_o;
  (* KEEP="TRUE" *) wire n9272_o;
  (* KEEP="TRUE" *) wire n9273_o;
  (* KEEP="TRUE" *) wire n9275_o;
  (* KEEP="TRUE" *) wire n9276_o;
  (* KEEP="TRUE" *) wire n9277_o;
  (* KEEP="TRUE" *) wire n9279_o;
  (* KEEP="TRUE" *) wire n9280_o;
  (* KEEP="TRUE" *) wire n9282_o;
  (* KEEP="TRUE" *) wire n9283_o;
  (* KEEP="TRUE" *) wire n9284_o;
  (* KEEP="TRUE" *) wire n9286_o;
  (* KEEP="TRUE" *) wire n9290_o;
  (* KEEP="TRUE" *) wire n9291_o;
  (* KEEP="TRUE" *) wire n9293_o;
  (* KEEP="TRUE" *) wire n9294_o;
  (* KEEP="TRUE" *) wire n9295_o;
  (* KEEP="TRUE" *) wire n9297_o;
  (* KEEP="TRUE" *) wire n9298_o;
  (* KEEP="TRUE" *) wire n9300_o;
  (* KEEP="TRUE" *) wire n9301_o;
  (* KEEP="TRUE" *) wire n9302_o;
  (* KEEP="TRUE" *) wire n9304_o;
  (* KEEP="TRUE" *) wire n9308_o;
  (* KEEP="TRUE" *) wire n9309_o;
  (* KEEP="TRUE" *) wire n9311_o;
  (* KEEP="TRUE" *) wire n9312_o;
  (* KEEP="TRUE" *) wire n9313_o;
  (* KEEP="TRUE" *) wire n9315_o;
  (* KEEP="TRUE" *) wire n9316_o;
  (* KEEP="TRUE" *) wire n9318_o;
  (* KEEP="TRUE" *) wire n9319_o;
  (* KEEP="TRUE" *) wire n9320_o;
  (* KEEP="TRUE" *) wire n9322_o;
  (* KEEP="TRUE" *) wire n9326_o;
  (* KEEP="TRUE" *) wire n9327_o;
  (* KEEP="TRUE" *) wire n9329_o;
  (* KEEP="TRUE" *) wire n9330_o;
  (* KEEP="TRUE" *) wire n9331_o;
  (* KEEP="TRUE" *) wire n9333_o;
  (* KEEP="TRUE" *) wire n9334_o;
  (* KEEP="TRUE" *) wire n9336_o;
  (* KEEP="TRUE" *) wire n9337_o;
  (* KEEP="TRUE" *) wire n9338_o;
  (* KEEP="TRUE" *) wire n9340_o;
  (* KEEP="TRUE" *) wire n9344_o;
  (* KEEP="TRUE" *) wire n9345_o;
  (* KEEP="TRUE" *) wire n9347_o;
  (* KEEP="TRUE" *) wire n9348_o;
  (* KEEP="TRUE" *) wire n9349_o;
  (* KEEP="TRUE" *) wire n9351_o;
  (* KEEP="TRUE" *) wire n9352_o;
  (* KEEP="TRUE" *) wire n9354_o;
  (* KEEP="TRUE" *) wire n9355_o;
  (* KEEP="TRUE" *) wire n9356_o;
  (* KEEP="TRUE" *) wire n9358_o;
  (* KEEP="TRUE" *) wire n9362_o;
  (* KEEP="TRUE" *) wire n9363_o;
  (* KEEP="TRUE" *) wire n9365_o;
  (* KEEP="TRUE" *) wire n9366_o;
  (* KEEP="TRUE" *) wire n9367_o;
  (* KEEP="TRUE" *) wire n9369_o;
  (* KEEP="TRUE" *) wire n9370_o;
  (* KEEP="TRUE" *) wire n9372_o;
  (* KEEP="TRUE" *) wire n9373_o;
  (* KEEP="TRUE" *) wire n9374_o;
  (* KEEP="TRUE" *) wire n9376_o;
  (* KEEP="TRUE" *) wire n9380_o;
  (* KEEP="TRUE" *) wire n9381_o;
  (* KEEP="TRUE" *) wire n9383_o;
  (* KEEP="TRUE" *) wire n9384_o;
  (* KEEP="TRUE" *) wire n9385_o;
  (* KEEP="TRUE" *) wire n9387_o;
  (* KEEP="TRUE" *) wire n9388_o;
  (* KEEP="TRUE" *) wire n9390_o;
  (* KEEP="TRUE" *) wire n9391_o;
  (* KEEP="TRUE" *) wire n9392_o;
  (* KEEP="TRUE" *) wire n9394_o;
  (* KEEP="TRUE" *) wire n9398_o;
  (* KEEP="TRUE" *) wire n9399_o;
  (* KEEP="TRUE" *) wire n9401_o;
  (* KEEP="TRUE" *) wire n9402_o;
  (* KEEP="TRUE" *) wire n9403_o;
  (* KEEP="TRUE" *) wire n9405_o;
  (* KEEP="TRUE" *) wire n9406_o;
  (* KEEP="TRUE" *) wire n9408_o;
  (* KEEP="TRUE" *) wire n9409_o;
  (* KEEP="TRUE" *) wire n9410_o;
  (* KEEP="TRUE" *) wire n9412_o;
  (* KEEP="TRUE" *) wire n9416_o;
  (* KEEP="TRUE" *) wire n9417_o;
  (* KEEP="TRUE" *) wire n9419_o;
  (* KEEP="TRUE" *) wire n9420_o;
  (* KEEP="TRUE" *) wire n9421_o;
  (* KEEP="TRUE" *) wire n9423_o;
  (* KEEP="TRUE" *) wire n9424_o;
  (* KEEP="TRUE" *) wire n9426_o;
  (* KEEP="TRUE" *) wire n9427_o;
  (* KEEP="TRUE" *) wire n9428_o;
  (* KEEP="TRUE" *) wire n9430_o;
  (* KEEP="TRUE" *) wire n9434_o;
  (* KEEP="TRUE" *) wire n9435_o;
  (* KEEP="TRUE" *) wire n9437_o;
  (* KEEP="TRUE" *) wire n9438_o;
  (* KEEP="TRUE" *) wire n9439_o;
  (* KEEP="TRUE" *) wire n9441_o;
  (* KEEP="TRUE" *) wire n9442_o;
  (* KEEP="TRUE" *) wire n9444_o;
  (* KEEP="TRUE" *) wire n9445_o;
  (* KEEP="TRUE" *) wire n9446_o;
  (* KEEP="TRUE" *) wire n9448_o;
  (* KEEP="TRUE" *) wire n9452_o;
  (* KEEP="TRUE" *) wire n9453_o;
  (* KEEP="TRUE" *) wire n9455_o;
  (* KEEP="TRUE" *) wire n9456_o;
  (* KEEP="TRUE" *) wire n9457_o;
  (* KEEP="TRUE" *) wire n9459_o;
  (* KEEP="TRUE" *) wire n9460_o;
  (* KEEP="TRUE" *) wire n9462_o;
  (* KEEP="TRUE" *) wire n9463_o;
  (* KEEP="TRUE" *) wire n9464_o;
  (* KEEP="TRUE" *) wire n9466_o;
  (* KEEP="TRUE" *) wire n9470_o;
  (* KEEP="TRUE" *) wire n9471_o;
  (* KEEP="TRUE" *) wire n9473_o;
  (* KEEP="TRUE" *) wire n9474_o;
  (* KEEP="TRUE" *) wire n9475_o;
  (* KEEP="TRUE" *) wire n9477_o;
  (* KEEP="TRUE" *) wire n9478_o;
  (* KEEP="TRUE" *) wire n9480_o;
  (* KEEP="TRUE" *) wire n9481_o;
  (* KEEP="TRUE" *) wire n9482_o;
  (* KEEP="TRUE" *) wire n9484_o;
  (* KEEP="TRUE" *) wire n9488_o;
  (* KEEP="TRUE" *) wire n9489_o;
  (* KEEP="TRUE" *) wire n9491_o;
  (* KEEP="TRUE" *) wire n9492_o;
  (* KEEP="TRUE" *) wire n9493_o;
  (* KEEP="TRUE" *) wire n9495_o;
  (* KEEP="TRUE" *) wire n9496_o;
  (* KEEP="TRUE" *) wire n9498_o;
  (* KEEP="TRUE" *) wire n9499_o;
  (* KEEP="TRUE" *) wire n9500_o;
  (* KEEP="TRUE" *) wire n9502_o;
  (* KEEP="TRUE" *) wire n9506_o;
  (* KEEP="TRUE" *) wire n9507_o;
  (* KEEP="TRUE" *) wire n9509_o;
  (* KEEP="TRUE" *) wire n9510_o;
  (* KEEP="TRUE" *) wire n9511_o;
  (* KEEP="TRUE" *) wire n9513_o;
  (* KEEP="TRUE" *) wire n9514_o;
  (* KEEP="TRUE" *) wire n9516_o;
  (* KEEP="TRUE" *) wire n9517_o;
  (* KEEP="TRUE" *) wire n9518_o;
  (* KEEP="TRUE" *) wire n9520_o;
  (* KEEP="TRUE" *) wire n9524_o;
  (* KEEP="TRUE" *) wire n9525_o;
  (* KEEP="TRUE" *) wire n9527_o;
  (* KEEP="TRUE" *) wire n9528_o;
  (* KEEP="TRUE" *) wire n9529_o;
  (* KEEP="TRUE" *) wire n9531_o;
  (* KEEP="TRUE" *) wire n9532_o;
  (* KEEP="TRUE" *) wire n9534_o;
  (* KEEP="TRUE" *) wire n9535_o;
  (* KEEP="TRUE" *) wire n9536_o;
  (* KEEP="TRUE" *) wire n9538_o;
  (* KEEP="TRUE" *) wire n9542_o;
  (* KEEP="TRUE" *) wire n9543_o;
  (* KEEP="TRUE" *) wire n9545_o;
  (* KEEP="TRUE" *) wire n9546_o;
  (* KEEP="TRUE" *) wire n9547_o;
  (* KEEP="TRUE" *) wire n9549_o;
  (* KEEP="TRUE" *) wire n9550_o;
  (* KEEP="TRUE" *) wire n9552_o;
  (* KEEP="TRUE" *) wire n9553_o;
  (* KEEP="TRUE" *) wire n9554_o;
  (* KEEP="TRUE" *) wire n9556_o;
  (* KEEP="TRUE" *) wire n9560_o;
  (* KEEP="TRUE" *) wire n9561_o;
  (* KEEP="TRUE" *) wire n9563_o;
  (* KEEP="TRUE" *) wire n9564_o;
  (* KEEP="TRUE" *) wire n9565_o;
  (* KEEP="TRUE" *) wire n9567_o;
  (* KEEP="TRUE" *) wire n9568_o;
  (* KEEP="TRUE" *) wire n9570_o;
  (* KEEP="TRUE" *) wire n9571_o;
  (* KEEP="TRUE" *) wire n9572_o;
  (* KEEP="TRUE" *) wire n9574_o;
  (* KEEP="TRUE" *) wire n9578_o;
  (* KEEP="TRUE" *) wire n9579_o;
  (* KEEP="TRUE" *) wire n9581_o;
  (* KEEP="TRUE" *) wire n9582_o;
  (* KEEP="TRUE" *) wire n9583_o;
  (* KEEP="TRUE" *) wire n9585_o;
  (* KEEP="TRUE" *) wire n9586_o;
  (* KEEP="TRUE" *) wire n9588_o;
  (* KEEP="TRUE" *) wire n9589_o;
  (* KEEP="TRUE" *) wire n9590_o;
  (* KEEP="TRUE" *) wire n9592_o;
  (* KEEP="TRUE" *) wire n9596_o;
  (* KEEP="TRUE" *) wire n9597_o;
  (* KEEP="TRUE" *) wire n9599_o;
  (* KEEP="TRUE" *) wire n9600_o;
  (* KEEP="TRUE" *) wire n9601_o;
  (* KEEP="TRUE" *) wire n9603_o;
  (* KEEP="TRUE" *) wire n9604_o;
  (* KEEP="TRUE" *) wire n9606_o;
  (* KEEP="TRUE" *) wire n9607_o;
  (* KEEP="TRUE" *) wire n9608_o;
  (* KEEP="TRUE" *) wire n9610_o;
  (* KEEP="TRUE" *) wire n9614_o;
  (* KEEP="TRUE" *) wire n9615_o;
  (* KEEP="TRUE" *) wire n9617_o;
  (* KEEP="TRUE" *) wire n9618_o;
  (* KEEP="TRUE" *) wire n9619_o;
  (* KEEP="TRUE" *) wire n9621_o;
  (* KEEP="TRUE" *) wire n9622_o;
  (* KEEP="TRUE" *) wire n9624_o;
  (* KEEP="TRUE" *) wire n9625_o;
  (* KEEP="TRUE" *) wire n9626_o;
  (* KEEP="TRUE" *) wire n9628_o;
  (* KEEP="TRUE" *) wire n9632_o;
  (* KEEP="TRUE" *) wire n9633_o;
  (* KEEP="TRUE" *) wire n9635_o;
  (* KEEP="TRUE" *) wire n9636_o;
  (* KEEP="TRUE" *) wire n9637_o;
  (* KEEP="TRUE" *) wire n9639_o;
  (* KEEP="TRUE" *) wire n9640_o;
  (* KEEP="TRUE" *) wire n9642_o;
  (* KEEP="TRUE" *) wire n9643_o;
  (* KEEP="TRUE" *) wire n9644_o;
  (* KEEP="TRUE" *) wire n9646_o;
  (* KEEP="TRUE" *) wire n9650_o;
  (* KEEP="TRUE" *) wire n9651_o;
  (* KEEP="TRUE" *) wire n9653_o;
  (* KEEP="TRUE" *) wire n9654_o;
  (* KEEP="TRUE" *) wire n9655_o;
  (* KEEP="TRUE" *) wire n9657_o;
  (* KEEP="TRUE" *) wire n9658_o;
  (* KEEP="TRUE" *) wire n9660_o;
  (* KEEP="TRUE" *) wire n9661_o;
  (* KEEP="TRUE" *) wire n9662_o;
  (* KEEP="TRUE" *) wire n9664_o;
  (* KEEP="TRUE" *) wire n9668_o;
  (* KEEP="TRUE" *) wire n9669_o;
  (* KEEP="TRUE" *) wire n9671_o;
  (* KEEP="TRUE" *) wire n9672_o;
  (* KEEP="TRUE" *) wire n9673_o;
  (* KEEP="TRUE" *) wire n9675_o;
  (* KEEP="TRUE" *) wire n9676_o;
  (* KEEP="TRUE" *) wire n9678_o;
  (* KEEP="TRUE" *) wire n9679_o;
  (* KEEP="TRUE" *) wire n9680_o;
  (* KEEP="TRUE" *) wire n9682_o;
  (* KEEP="TRUE" *) wire n9686_o;
  (* KEEP="TRUE" *) wire n9687_o;
  (* KEEP="TRUE" *) wire n9689_o;
  (* KEEP="TRUE" *) wire n9690_o;
  (* KEEP="TRUE" *) wire n9691_o;
  (* KEEP="TRUE" *) wire n9693_o;
  (* KEEP="TRUE" *) wire n9694_o;
  (* KEEP="TRUE" *) wire n9696_o;
  (* KEEP="TRUE" *) wire n9697_o;
  (* KEEP="TRUE" *) wire n9698_o;
  (* KEEP="TRUE" *) wire n9700_o;
  (* KEEP="TRUE" *) wire n9704_o;
  (* KEEP="TRUE" *) wire n9705_o;
  (* KEEP="TRUE" *) wire n9707_o;
  (* KEEP="TRUE" *) wire n9708_o;
  (* KEEP="TRUE" *) wire n9709_o;
  (* KEEP="TRUE" *) wire n9711_o;
  (* KEEP="TRUE" *) wire n9712_o;
  (* KEEP="TRUE" *) wire n9714_o;
  (* KEEP="TRUE" *) wire n9715_o;
  (* KEEP="TRUE" *) wire n9716_o;
  (* KEEP="TRUE" *) wire n9718_o;
  (* KEEP="TRUE" *) wire n9722_o;
  (* KEEP="TRUE" *) wire n9723_o;
  (* KEEP="TRUE" *) wire n9725_o;
  (* KEEP="TRUE" *) wire n9726_o;
  (* KEEP="TRUE" *) wire n9727_o;
  (* KEEP="TRUE" *) wire n9729_o;
  (* KEEP="TRUE" *) wire n9730_o;
  (* KEEP="TRUE" *) wire n9732_o;
  (* KEEP="TRUE" *) wire n9733_o;
  (* KEEP="TRUE" *) wire n9734_o;
  (* KEEP="TRUE" *) wire n9736_o;
  (* KEEP="TRUE" *) wire n9740_o;
  (* KEEP="TRUE" *) wire n9741_o;
  (* KEEP="TRUE" *) wire n9743_o;
  (* KEEP="TRUE" *) wire n9744_o;
  (* KEEP="TRUE" *) wire n9745_o;
  (* KEEP="TRUE" *) wire n9747_o;
  (* KEEP="TRUE" *) wire n9748_o;
  (* KEEP="TRUE" *) wire n9750_o;
  (* KEEP="TRUE" *) wire n9751_o;
  (* KEEP="TRUE" *) wire n9752_o;
  (* KEEP="TRUE" *) wire n9754_o;
  (* KEEP="TRUE" *) wire n9758_o;
  (* KEEP="TRUE" *) wire n9759_o;
  (* KEEP="TRUE" *) wire n9761_o;
  (* KEEP="TRUE" *) wire n9762_o;
  (* KEEP="TRUE" *) wire n9763_o;
  (* KEEP="TRUE" *) wire n9765_o;
  (* KEEP="TRUE" *) wire n9766_o;
  (* KEEP="TRUE" *) wire n9768_o;
  (* KEEP="TRUE" *) wire n9769_o;
  (* KEEP="TRUE" *) wire n9770_o;
  (* KEEP="TRUE" *) wire n9772_o;
  (* KEEP="TRUE" *) wire n9776_o;
  (* KEEP="TRUE" *) wire n9777_o;
  (* KEEP="TRUE" *) wire n9779_o;
  (* KEEP="TRUE" *) wire n9780_o;
  (* KEEP="TRUE" *) wire n9781_o;
  (* KEEP="TRUE" *) wire n9783_o;
  (* KEEP="TRUE" *) wire n9784_o;
  (* KEEP="TRUE" *) wire n9786_o;
  (* KEEP="TRUE" *) wire n9787_o;
  (* KEEP="TRUE" *) wire n9788_o;
  (* KEEP="TRUE" *) wire n9790_o;
  (* KEEP="TRUE" *) wire n9794_o;
  (* KEEP="TRUE" *) wire n9795_o;
  (* KEEP="TRUE" *) wire n9797_o;
  (* KEEP="TRUE" *) wire n9798_o;
  (* KEEP="TRUE" *) wire n9799_o;
  (* KEEP="TRUE" *) wire n9801_o;
  (* KEEP="TRUE" *) wire n9802_o;
  (* KEEP="TRUE" *) wire n9804_o;
  (* KEEP="TRUE" *) wire n9805_o;
  (* KEEP="TRUE" *) wire n9806_o;
  (* KEEP="TRUE" *) wire n9808_o;
  (* KEEP="TRUE" *) wire n9812_o;
  (* KEEP="TRUE" *) wire n9813_o;
  (* KEEP="TRUE" *) wire n9815_o;
  (* KEEP="TRUE" *) wire n9816_o;
  (* KEEP="TRUE" *) wire n9817_o;
  (* KEEP="TRUE" *) wire n9819_o;
  (* KEEP="TRUE" *) wire n9820_o;
  (* KEEP="TRUE" *) wire n9822_o;
  (* KEEP="TRUE" *) wire n9823_o;
  (* KEEP="TRUE" *) wire n9824_o;
  (* KEEP="TRUE" *) wire n9826_o;
  (* KEEP="TRUE" *) wire n9830_o;
  (* KEEP="TRUE" *) wire n9831_o;
  (* KEEP="TRUE" *) wire n9833_o;
  (* KEEP="TRUE" *) wire n9834_o;
  (* KEEP="TRUE" *) wire n9835_o;
  (* KEEP="TRUE" *) wire n9837_o;
  (* KEEP="TRUE" *) wire n9838_o;
  (* KEEP="TRUE" *) wire n9840_o;
  (* KEEP="TRUE" *) wire n9841_o;
  (* KEEP="TRUE" *) wire n9842_o;
  (* KEEP="TRUE" *) wire n9844_o;
  (* KEEP="TRUE" *) wire n9848_o;
  (* KEEP="TRUE" *) wire n9849_o;
  (* KEEP="TRUE" *) wire n9851_o;
  (* KEEP="TRUE" *) wire n9852_o;
  (* KEEP="TRUE" *) wire n9853_o;
  (* KEEP="TRUE" *) wire n9855_o;
  (* KEEP="TRUE" *) wire n9856_o;
  (* KEEP="TRUE" *) wire n9858_o;
  (* KEEP="TRUE" *) wire n9859_o;
  (* KEEP="TRUE" *) wire n9860_o;
  (* KEEP="TRUE" *) wire n9862_o;
  (* KEEP="TRUE" *) wire n9866_o;
  (* KEEP="TRUE" *) wire n9867_o;
  (* KEEP="TRUE" *) wire n9869_o;
  (* KEEP="TRUE" *) wire n9870_o;
  (* KEEP="TRUE" *) wire n9871_o;
  (* KEEP="TRUE" *) wire n9873_o;
  (* KEEP="TRUE" *) wire n9874_o;
  (* KEEP="TRUE" *) wire n9876_o;
  (* KEEP="TRUE" *) wire n9877_o;
  (* KEEP="TRUE" *) wire n9878_o;
  (* KEEP="TRUE" *) wire n9880_o;
  (* KEEP="TRUE" *) wire n9884_o;
  (* KEEP="TRUE" *) wire n9885_o;
  (* KEEP="TRUE" *) wire n9887_o;
  (* KEEP="TRUE" *) wire n9888_o;
  (* KEEP="TRUE" *) wire n9889_o;
  (* KEEP="TRUE" *) wire n9891_o;
  (* KEEP="TRUE" *) wire n9892_o;
  (* KEEP="TRUE" *) wire n9894_o;
  (* KEEP="TRUE" *) wire n9895_o;
  (* KEEP="TRUE" *) wire n9896_o;
  (* KEEP="TRUE" *) wire n9898_o;
  (* KEEP="TRUE" *) wire n9902_o;
  (* KEEP="TRUE" *) wire n9903_o;
  (* KEEP="TRUE" *) wire n9905_o;
  (* KEEP="TRUE" *) wire n9906_o;
  (* KEEP="TRUE" *) wire n9907_o;
  (* KEEP="TRUE" *) wire n9909_o;
  (* KEEP="TRUE" *) wire n9910_o;
  (* KEEP="TRUE" *) wire n9912_o;
  (* KEEP="TRUE" *) wire n9913_o;
  (* KEEP="TRUE" *) wire n9914_o;
  (* KEEP="TRUE" *) wire n9916_o;
  (* KEEP="TRUE" *) wire n9920_o;
  (* KEEP="TRUE" *) wire n9921_o;
  (* KEEP="TRUE" *) wire n9923_o;
  (* KEEP="TRUE" *) wire n9924_o;
  (* KEEP="TRUE" *) wire n9925_o;
  (* KEEP="TRUE" *) wire n9927_o;
  (* KEEP="TRUE" *) wire n9928_o;
  (* KEEP="TRUE" *) wire n9930_o;
  (* KEEP="TRUE" *) wire n9931_o;
  (* KEEP="TRUE" *) wire n9932_o;
  (* KEEP="TRUE" *) wire n9934_o;
  (* KEEP="TRUE" *) wire n9938_o;
  (* KEEP="TRUE" *) wire n9939_o;
  (* KEEP="TRUE" *) wire n9941_o;
  (* KEEP="TRUE" *) wire n9942_o;
  (* KEEP="TRUE" *) wire n9943_o;
  (* KEEP="TRUE" *) wire n9945_o;
  (* KEEP="TRUE" *) wire n9946_o;
  (* KEEP="TRUE" *) wire n9948_o;
  (* KEEP="TRUE" *) wire n9949_o;
  (* KEEP="TRUE" *) wire n9950_o;
  (* KEEP="TRUE" *) wire n9952_o;
  (* KEEP="TRUE" *) wire n9956_o;
  (* KEEP="TRUE" *) wire n9957_o;
  (* KEEP="TRUE" *) wire n9959_o;
  (* KEEP="TRUE" *) wire n9960_o;
  (* KEEP="TRUE" *) wire n9961_o;
  (* KEEP="TRUE" *) wire n9963_o;
  (* KEEP="TRUE" *) wire n9964_o;
  (* KEEP="TRUE" *) wire n9966_o;
  (* KEEP="TRUE" *) wire n9967_o;
  (* KEEP="TRUE" *) wire n9968_o;
  (* KEEP="TRUE" *) wire n9970_o;
  (* KEEP="TRUE" *) wire n9974_o;
  (* KEEP="TRUE" *) wire n9975_o;
  (* KEEP="TRUE" *) wire n9977_o;
  (* KEEP="TRUE" *) wire n9978_o;
  (* KEEP="TRUE" *) wire n9979_o;
  (* KEEP="TRUE" *) wire n9981_o;
  (* KEEP="TRUE" *) wire n9982_o;
  (* KEEP="TRUE" *) wire n9984_o;
  (* KEEP="TRUE" *) wire n9985_o;
  (* KEEP="TRUE" *) wire n9986_o;
  (* KEEP="TRUE" *) wire n9988_o;
  (* KEEP="TRUE" *) wire n9992_o;
  (* KEEP="TRUE" *) wire n9993_o;
  (* KEEP="TRUE" *) wire n9995_o;
  (* KEEP="TRUE" *) wire n9996_o;
  (* KEEP="TRUE" *) wire n9997_o;
  (* KEEP="TRUE" *) wire n9999_o;
  (* KEEP="TRUE" *) wire n10000_o;
  (* KEEP="TRUE" *) wire n10002_o;
  (* KEEP="TRUE" *) wire n10003_o;
  (* KEEP="TRUE" *) wire n10004_o;
  (* KEEP="TRUE" *) wire n10006_o;
  (* KEEP="TRUE" *) wire n10010_o;
  (* KEEP="TRUE" *) wire n10011_o;
  (* KEEP="TRUE" *) wire n10013_o;
  (* KEEP="TRUE" *) wire n10014_o;
  (* KEEP="TRUE" *) wire n10015_o;
  (* KEEP="TRUE" *) wire n10017_o;
  (* KEEP="TRUE" *) wire n10018_o;
  (* KEEP="TRUE" *) wire n10020_o;
  (* KEEP="TRUE" *) wire n10021_o;
  (* KEEP="TRUE" *) wire n10022_o;
  (* KEEP="TRUE" *) wire n10024_o;
  (* KEEP="TRUE" *) wire n10028_o;
  (* KEEP="TRUE" *) wire n10029_o;
  (* KEEP="TRUE" *) wire n10031_o;
  (* KEEP="TRUE" *) wire n10032_o;
  (* KEEP="TRUE" *) wire n10033_o;
  (* KEEP="TRUE" *) wire n10035_o;
  (* KEEP="TRUE" *) wire n10036_o;
  (* KEEP="TRUE" *) wire n10038_o;
  (* KEEP="TRUE" *) wire n10039_o;
  (* KEEP="TRUE" *) wire n10040_o;
  (* KEEP="TRUE" *) wire n10042_o;
  (* KEEP="TRUE" *) wire n10046_o;
  (* KEEP="TRUE" *) wire n10047_o;
  (* KEEP="TRUE" *) wire n10049_o;
  (* KEEP="TRUE" *) wire n10050_o;
  (* KEEP="TRUE" *) wire n10051_o;
  (* KEEP="TRUE" *) wire n10053_o;
  (* KEEP="TRUE" *) wire n10054_o;
  (* KEEP="TRUE" *) wire n10056_o;
  (* KEEP="TRUE" *) wire n10057_o;
  (* KEEP="TRUE" *) wire n10058_o;
  (* KEEP="TRUE" *) wire n10060_o;
  (* KEEP="TRUE" *) wire n10064_o;
  (* KEEP="TRUE" *) wire n10065_o;
  (* KEEP="TRUE" *) wire n10067_o;
  (* KEEP="TRUE" *) wire n10068_o;
  (* KEEP="TRUE" *) wire n10069_o;
  (* KEEP="TRUE" *) wire n10071_o;
  (* KEEP="TRUE" *) wire n10072_o;
  (* KEEP="TRUE" *) wire n10074_o;
  (* KEEP="TRUE" *) wire n10075_o;
  (* KEEP="TRUE" *) wire n10076_o;
  (* KEEP="TRUE" *) wire n10078_o;
  (* KEEP="TRUE" *) wire n10082_o;
  (* KEEP="TRUE" *) wire n10083_o;
  (* KEEP="TRUE" *) wire n10085_o;
  (* KEEP="TRUE" *) wire n10086_o;
  (* KEEP="TRUE" *) wire n10087_o;
  (* KEEP="TRUE" *) wire n10089_o;
  (* KEEP="TRUE" *) wire n10090_o;
  (* KEEP="TRUE" *) wire n10092_o;
  (* KEEP="TRUE" *) wire n10093_o;
  (* KEEP="TRUE" *) wire n10094_o;
  (* KEEP="TRUE" *) wire n10096_o;
  (* KEEP="TRUE" *) wire n10100_o;
  (* KEEP="TRUE" *) wire n10101_o;
  (* KEEP="TRUE" *) wire n10103_o;
  (* KEEP="TRUE" *) wire n10104_o;
  (* KEEP="TRUE" *) wire n10105_o;
  (* KEEP="TRUE" *) wire n10107_o;
  (* KEEP="TRUE" *) wire n10108_o;
  (* KEEP="TRUE" *) wire n10110_o;
  (* KEEP="TRUE" *) wire n10111_o;
  (* KEEP="TRUE" *) wire n10112_o;
  (* KEEP="TRUE" *) wire n10114_o;
  (* KEEP="TRUE" *) wire n10118_o;
  (* KEEP="TRUE" *) wire n10119_o;
  (* KEEP="TRUE" *) wire n10121_o;
  (* KEEP="TRUE" *) wire n10122_o;
  (* KEEP="TRUE" *) wire n10123_o;
  (* KEEP="TRUE" *) wire n10125_o;
  (* KEEP="TRUE" *) wire n10126_o;
  (* KEEP="TRUE" *) wire n10128_o;
  (* KEEP="TRUE" *) wire n10129_o;
  (* KEEP="TRUE" *) wire n10130_o;
  (* KEEP="TRUE" *) wire n10132_o;
  (* KEEP="TRUE" *) wire n10136_o;
  (* KEEP="TRUE" *) wire n10137_o;
  (* KEEP="TRUE" *) wire n10139_o;
  (* KEEP="TRUE" *) wire n10140_o;
  (* KEEP="TRUE" *) wire n10141_o;
  (* KEEP="TRUE" *) wire n10143_o;
  (* KEEP="TRUE" *) wire n10144_o;
  (* KEEP="TRUE" *) wire n10146_o;
  (* KEEP="TRUE" *) wire n10147_o;
  (* KEEP="TRUE" *) wire n10148_o;
  (* KEEP="TRUE" *) wire n10150_o;
  (* KEEP="TRUE" *) wire n10154_o;
  (* KEEP="TRUE" *) wire n10155_o;
  (* KEEP="TRUE" *) wire n10157_o;
  (* KEEP="TRUE" *) wire n10158_o;
  (* KEEP="TRUE" *) wire n10159_o;
  (* KEEP="TRUE" *) wire n10161_o;
  (* KEEP="TRUE" *) wire n10162_o;
  (* KEEP="TRUE" *) wire n10164_o;
  (* KEEP="TRUE" *) wire n10165_o;
  (* KEEP="TRUE" *) wire n10166_o;
  (* KEEP="TRUE" *) wire n10168_o;
  (* KEEP="TRUE" *) wire n10172_o;
  (* KEEP="TRUE" *) wire n10173_o;
  (* KEEP="TRUE" *) wire n10175_o;
  (* KEEP="TRUE" *) wire n10176_o;
  (* KEEP="TRUE" *) wire n10177_o;
  (* KEEP="TRUE" *) wire n10179_o;
  (* KEEP="TRUE" *) wire n10180_o;
  (* KEEP="TRUE" *) wire n10182_o;
  (* KEEP="TRUE" *) wire n10183_o;
  (* KEEP="TRUE" *) wire n10184_o;
  (* KEEP="TRUE" *) wire n10186_o;
  (* KEEP="TRUE" *) wire n10190_o;
  (* KEEP="TRUE" *) wire n10191_o;
  (* KEEP="TRUE" *) wire n10193_o;
  (* KEEP="TRUE" *) wire n10194_o;
  (* KEEP="TRUE" *) wire n10195_o;
  (* KEEP="TRUE" *) wire n10197_o;
  (* KEEP="TRUE" *) wire n10198_o;
  (* KEEP="TRUE" *) wire n10200_o;
  (* KEEP="TRUE" *) wire n10201_o;
  (* KEEP="TRUE" *) wire n10202_o;
  (* KEEP="TRUE" *) wire n10204_o;
  (* KEEP="TRUE" *) wire n10208_o;
  (* KEEP="TRUE" *) wire n10209_o;
  (* KEEP="TRUE" *) wire n10211_o;
  (* KEEP="TRUE" *) wire n10212_o;
  (* KEEP="TRUE" *) wire n10213_o;
  (* KEEP="TRUE" *) wire n10215_o;
  (* KEEP="TRUE" *) wire n10216_o;
  (* KEEP="TRUE" *) wire n10218_o;
  (* KEEP="TRUE" *) wire n10219_o;
  (* KEEP="TRUE" *) wire n10220_o;
  (* KEEP="TRUE" *) wire n10222_o;
  (* KEEP="TRUE" *) wire n10226_o;
  (* KEEP="TRUE" *) wire n10227_o;
  (* KEEP="TRUE" *) wire n10229_o;
  (* KEEP="TRUE" *) wire n10230_o;
  (* KEEP="TRUE" *) wire n10231_o;
  (* KEEP="TRUE" *) wire n10233_o;
  (* KEEP="TRUE" *) wire n10234_o;
  (* KEEP="TRUE" *) wire n10236_o;
  (* KEEP="TRUE" *) wire n10237_o;
  (* KEEP="TRUE" *) wire n10238_o;
  (* KEEP="TRUE" *) wire n10240_o;
  (* KEEP="TRUE" *) wire n10244_o;
  (* KEEP="TRUE" *) wire n10245_o;
  (* KEEP="TRUE" *) wire n10247_o;
  (* KEEP="TRUE" *) wire n10248_o;
  (* KEEP="TRUE" *) wire n10249_o;
  (* KEEP="TRUE" *) wire n10251_o;
  (* KEEP="TRUE" *) wire n10252_o;
  (* KEEP="TRUE" *) wire n10254_o;
  (* KEEP="TRUE" *) wire n10255_o;
  (* KEEP="TRUE" *) wire n10256_o;
  (* KEEP="TRUE" *) wire n10258_o;
  (* KEEP="TRUE" *) wire n10262_o;
  (* KEEP="TRUE" *) wire n10263_o;
  (* KEEP="TRUE" *) wire n10265_o;
  (* KEEP="TRUE" *) wire n10266_o;
  (* KEEP="TRUE" *) wire n10267_o;
  (* KEEP="TRUE" *) wire n10269_o;
  (* KEEP="TRUE" *) wire n10270_o;
  (* KEEP="TRUE" *) wire n10272_o;
  (* KEEP="TRUE" *) wire n10273_o;
  (* KEEP="TRUE" *) wire n10274_o;
  (* KEEP="TRUE" *) wire n10276_o;
  (* KEEP="TRUE" *) wire n10280_o;
  (* KEEP="TRUE" *) wire n10281_o;
  (* KEEP="TRUE" *) wire n10283_o;
  (* KEEP="TRUE" *) wire n10284_o;
  (* KEEP="TRUE" *) wire n10285_o;
  (* KEEP="TRUE" *) wire n10287_o;
  (* KEEP="TRUE" *) wire n10288_o;
  (* KEEP="TRUE" *) wire n10290_o;
  (* KEEP="TRUE" *) wire n10291_o;
  (* KEEP="TRUE" *) wire n10292_o;
  (* KEEP="TRUE" *) wire n10294_o;
  (* KEEP="TRUE" *) wire n10298_o;
  (* KEEP="TRUE" *) wire n10299_o;
  (* KEEP="TRUE" *) wire n10301_o;
  (* KEEP="TRUE" *) wire n10302_o;
  (* KEEP="TRUE" *) wire n10303_o;
  (* KEEP="TRUE" *) wire n10305_o;
  (* KEEP="TRUE" *) wire n10306_o;
  (* KEEP="TRUE" *) wire n10308_o;
  (* KEEP="TRUE" *) wire n10309_o;
  (* KEEP="TRUE" *) wire n10310_o;
  (* KEEP="TRUE" *) wire n10312_o;
  (* KEEP="TRUE" *) wire n10316_o;
  (* KEEP="TRUE" *) wire n10317_o;
  (* KEEP="TRUE" *) wire n10319_o;
  (* KEEP="TRUE" *) wire n10320_o;
  (* KEEP="TRUE" *) wire n10321_o;
  (* KEEP="TRUE" *) wire n10323_o;
  (* KEEP="TRUE" *) wire n10324_o;
  (* KEEP="TRUE" *) wire n10326_o;
  (* KEEP="TRUE" *) wire n10327_o;
  (* KEEP="TRUE" *) wire n10328_o;
  (* KEEP="TRUE" *) wire n10330_o;
  (* KEEP="TRUE" *) wire n10334_o;
  (* KEEP="TRUE" *) wire n10335_o;
  (* KEEP="TRUE" *) wire n10337_o;
  (* KEEP="TRUE" *) wire n10338_o;
  (* KEEP="TRUE" *) wire n10339_o;
  (* KEEP="TRUE" *) wire n10341_o;
  (* KEEP="TRUE" *) wire n10342_o;
  (* KEEP="TRUE" *) wire n10344_o;
  (* KEEP="TRUE" *) wire n10345_o;
  (* KEEP="TRUE" *) wire n10346_o;
  (* KEEP="TRUE" *) wire n10348_o;
  (* KEEP="TRUE" *) wire n10352_o;
  (* KEEP="TRUE" *) wire n10353_o;
  (* KEEP="TRUE" *) wire n10355_o;
  (* KEEP="TRUE" *) wire n10356_o;
  (* KEEP="TRUE" *) wire n10357_o;
  (* KEEP="TRUE" *) wire n10359_o;
  (* KEEP="TRUE" *) wire n10360_o;
  (* KEEP="TRUE" *) wire n10362_o;
  (* KEEP="TRUE" *) wire n10363_o;
  (* KEEP="TRUE" *) wire n10364_o;
  (* KEEP="TRUE" *) wire n10366_o;
  (* KEEP="TRUE" *) wire n10370_o;
  (* KEEP="TRUE" *) wire n10371_o;
  (* KEEP="TRUE" *) wire n10373_o;
  (* KEEP="TRUE" *) wire n10374_o;
  (* KEEP="TRUE" *) wire n10375_o;
  (* KEEP="TRUE" *) wire n10377_o;
  (* KEEP="TRUE" *) wire n10378_o;
  (* KEEP="TRUE" *) wire n10380_o;
  (* KEEP="TRUE" *) wire n10381_o;
  (* KEEP="TRUE" *) wire n10382_o;
  (* KEEP="TRUE" *) wire n10384_o;
  (* KEEP="TRUE" *) wire n10388_o;
  (* KEEP="TRUE" *) wire n10389_o;
  (* KEEP="TRUE" *) wire n10391_o;
  (* KEEP="TRUE" *) wire n10392_o;
  (* KEEP="TRUE" *) wire n10393_o;
  (* KEEP="TRUE" *) wire n10395_o;
  (* KEEP="TRUE" *) wire n10396_o;
  (* KEEP="TRUE" *) wire n10398_o;
  (* KEEP="TRUE" *) wire n10399_o;
  (* KEEP="TRUE" *) wire n10400_o;
  (* KEEP="TRUE" *) wire n10402_o;
  (* KEEP="TRUE" *) wire n10406_o;
  (* KEEP="TRUE" *) wire n10407_o;
  (* KEEP="TRUE" *) wire n10409_o;
  (* KEEP="TRUE" *) wire n10410_o;
  (* KEEP="TRUE" *) wire n10411_o;
  (* KEEP="TRUE" *) wire n10413_o;
  (* KEEP="TRUE" *) wire n10414_o;
  (* KEEP="TRUE" *) wire n10416_o;
  (* KEEP="TRUE" *) wire n10417_o;
  (* KEEP="TRUE" *) wire n10418_o;
  (* KEEP="TRUE" *) wire n10420_o;
  (* KEEP="TRUE" *) wire n10424_o;
  (* KEEP="TRUE" *) wire n10425_o;
  (* KEEP="TRUE" *) wire n10427_o;
  (* KEEP="TRUE" *) wire n10428_o;
  (* KEEP="TRUE" *) wire n10429_o;
  (* KEEP="TRUE" *) wire n10431_o;
  (* KEEP="TRUE" *) wire n10432_o;
  (* KEEP="TRUE" *) wire n10434_o;
  (* KEEP="TRUE" *) wire n10435_o;
  (* KEEP="TRUE" *) wire n10436_o;
  (* KEEP="TRUE" *) wire n10438_o;
  (* KEEP="TRUE" *) wire n10442_o;
  (* KEEP="TRUE" *) wire n10443_o;
  (* KEEP="TRUE" *) wire n10445_o;
  (* KEEP="TRUE" *) wire n10446_o;
  (* KEEP="TRUE" *) wire n10447_o;
  (* KEEP="TRUE" *) wire n10449_o;
  (* KEEP="TRUE" *) wire n10450_o;
  (* KEEP="TRUE" *) wire n10452_o;
  (* KEEP="TRUE" *) wire n10453_o;
  (* KEEP="TRUE" *) wire n10454_o;
  (* KEEP="TRUE" *) wire n10456_o;
  (* KEEP="TRUE" *) wire n10460_o;
  (* KEEP="TRUE" *) wire n10461_o;
  (* KEEP="TRUE" *) wire n10463_o;
  (* KEEP="TRUE" *) wire n10464_o;
  (* KEEP="TRUE" *) wire n10465_o;
  (* KEEP="TRUE" *) wire n10467_o;
  (* KEEP="TRUE" *) wire n10468_o;
  (* KEEP="TRUE" *) wire n10470_o;
  (* KEEP="TRUE" *) wire n10471_o;
  (* KEEP="TRUE" *) wire n10472_o;
  (* KEEP="TRUE" *) wire n10474_o;
  (* KEEP="TRUE" *) wire n10478_o;
  (* KEEP="TRUE" *) wire n10479_o;
  (* KEEP="TRUE" *) wire n10481_o;
  (* KEEP="TRUE" *) wire n10482_o;
  (* KEEP="TRUE" *) wire n10483_o;
  (* KEEP="TRUE" *) wire n10485_o;
  (* KEEP="TRUE" *) wire n10486_o;
  (* KEEP="TRUE" *) wire n10488_o;
  (* KEEP="TRUE" *) wire n10489_o;
  (* KEEP="TRUE" *) wire n10490_o;
  (* KEEP="TRUE" *) wire n10492_o;
  (* KEEP="TRUE" *) wire n10497_o;
  (* KEEP="TRUE" *) wire n10499_o;
  (* KEEP="TRUE" *) wire n10501_o;
  (* KEEP="TRUE" *) wire n10503_o;
  (* KEEP="TRUE" *) wire n10505_o;
  (* KEEP="TRUE" *) wire n10507_o;
  (* KEEP="TRUE" *) wire [255:0] n10765_o;
  (* KEEP="TRUE" *) wire n10766_o;
  (* KEEP="TRUE" *) wire n10767_o;
  (* KEEP="TRUE" *) wire n10768_o;
  (* KEEP="TRUE" *) wire n10769_o;
  (* KEEP="TRUE" *) wire n10770_o;
  (* KEEP="TRUE" *) wire n10771_o;
  (* KEEP="TRUE" *) wire n10772_o;
  (* KEEP="TRUE" *) wire n10773_o;
  (* KEEP="TRUE" *) wire n10774_o;
  (* KEEP="TRUE" *) wire n10775_o;
  (* KEEP="TRUE" *) wire n10776_o;
  (* KEEP="TRUE" *) wire n10777_o;
  (* KEEP="TRUE" *) wire n10778_o;
  (* KEEP="TRUE" *) wire n10779_o;
  (* KEEP="TRUE" *) wire n10780_o;
  (* KEEP="TRUE" *) wire n10781_o;
  (* KEEP="TRUE" *) wire n10782_o;
  (* KEEP="TRUE" *) wire n10783_o;
  (* KEEP="TRUE" *) wire n10784_o;
  (* KEEP="TRUE" *) wire n10785_o;
  (* KEEP="TRUE" *) wire n10786_o;
  (* KEEP="TRUE" *) wire n10787_o;
  (* KEEP="TRUE" *) wire n10788_o;
  (* KEEP="TRUE" *) wire n10789_o;
  (* KEEP="TRUE" *) wire n10790_o;
  (* KEEP="TRUE" *) wire n10791_o;
  (* KEEP="TRUE" *) wire n10792_o;
  (* KEEP="TRUE" *) wire n10793_o;
  (* KEEP="TRUE" *) wire n10794_o;
  (* KEEP="TRUE" *) wire n10795_o;
  (* KEEP="TRUE" *) wire n10796_o;
  (* KEEP="TRUE" *) wire n10797_o;
  (* KEEP="TRUE" *) wire n10798_o;
  (* KEEP="TRUE" *) wire n10799_o;
  (* KEEP="TRUE" *) wire n10800_o;
  (* KEEP="TRUE" *) wire n10801_o;
  (* KEEP="TRUE" *) wire n10802_o;
  (* KEEP="TRUE" *) wire n10803_o;
  (* KEEP="TRUE" *) wire n10804_o;
  (* KEEP="TRUE" *) wire n10805_o;
  (* KEEP="TRUE" *) wire n10806_o;
  (* KEEP="TRUE" *) wire n10807_o;
  (* KEEP="TRUE" *) wire n10808_o;
  (* KEEP="TRUE" *) wire n10809_o;
  (* KEEP="TRUE" *) wire n10810_o;
  (* KEEP="TRUE" *) wire n10811_o;
  (* KEEP="TRUE" *) wire n10812_o;
  (* KEEP="TRUE" *) wire n10813_o;
  (* KEEP="TRUE" *) wire n10814_o;
  (* KEEP="TRUE" *) wire n10815_o;
  (* KEEP="TRUE" *) wire n10816_o;
  (* KEEP="TRUE" *) wire n10817_o;
  (* KEEP="TRUE" *) wire n10818_o;
  (* KEEP="TRUE" *) wire n10819_o;
  (* KEEP="TRUE" *) wire n10820_o;
  (* KEEP="TRUE" *) wire n10821_o;
  (* KEEP="TRUE" *) wire n10822_o;
  (* KEEP="TRUE" *) wire n10823_o;
  (* KEEP="TRUE" *) wire n10824_o;
  (* KEEP="TRUE" *) wire n10825_o;
  (* KEEP="TRUE" *) wire n10826_o;
  (* KEEP="TRUE" *) wire n10827_o;
  (* KEEP="TRUE" *) wire n10828_o;
  (* KEEP="TRUE" *) wire n10829_o;
  (* KEEP="TRUE" *) wire n10830_o;
  (* KEEP="TRUE" *) wire n10831_o;
  (* KEEP="TRUE" *) wire n10832_o;
  (* KEEP="TRUE" *) wire n10833_o;
  (* KEEP="TRUE" *) wire n10834_o;
  (* KEEP="TRUE" *) wire n10835_o;
  (* KEEP="TRUE" *) wire n10836_o;
  (* KEEP="TRUE" *) wire n10837_o;
  (* KEEP="TRUE" *) wire n10838_o;
  (* KEEP="TRUE" *) wire n10839_o;
  (* KEEP="TRUE" *) wire n10840_o;
  (* KEEP="TRUE" *) wire n10841_o;
  (* KEEP="TRUE" *) wire n10842_o;
  (* KEEP="TRUE" *) wire n10843_o;
  (* KEEP="TRUE" *) wire n10844_o;
  (* KEEP="TRUE" *) wire n10845_o;
  (* KEEP="TRUE" *) wire n10846_o;
  (* KEEP="TRUE" *) wire n10847_o;
  (* KEEP="TRUE" *) wire n10848_o;
  (* KEEP="TRUE" *) wire n10849_o;
  (* KEEP="TRUE" *) wire n10850_o;
  (* KEEP="TRUE" *) wire n10851_o;
  (* KEEP="TRUE" *) wire n10852_o;
  (* KEEP="TRUE" *) wire n10853_o;
  (* KEEP="TRUE" *) wire n10854_o;
  (* KEEP="TRUE" *) wire n10855_o;
  (* KEEP="TRUE" *) wire n10856_o;
  (* KEEP="TRUE" *) wire n10857_o;
  (* KEEP="TRUE" *) wire n10858_o;
  (* KEEP="TRUE" *) wire n10859_o;
  (* KEEP="TRUE" *) wire n10860_o;
  (* KEEP="TRUE" *) wire n10861_o;
  (* KEEP="TRUE" *) wire n10862_o;
  (* KEEP="TRUE" *) wire n10863_o;
  (* KEEP="TRUE" *) wire n10864_o;
  (* KEEP="TRUE" *) wire n10865_o;
  (* KEEP="TRUE" *) wire n10866_o;
  (* KEEP="TRUE" *) wire n10867_o;
  (* KEEP="TRUE" *) wire n10868_o;
  (* KEEP="TRUE" *) wire n10869_o;
  (* KEEP="TRUE" *) wire n10870_o;
  (* KEEP="TRUE" *) wire n10871_o;
  (* KEEP="TRUE" *) wire n10872_o;
  (* KEEP="TRUE" *) wire n10873_o;
  (* KEEP="TRUE" *) wire n10874_o;
  (* KEEP="TRUE" *) wire n10875_o;
  (* KEEP="TRUE" *) wire n10876_o;
  (* KEEP="TRUE" *) wire n10877_o;
  (* KEEP="TRUE" *) wire n10878_o;
  (* KEEP="TRUE" *) wire n10879_o;
  (* KEEP="TRUE" *) wire n10880_o;
  (* KEEP="TRUE" *) wire n10881_o;
  (* KEEP="TRUE" *) wire n10882_o;
  (* KEEP="TRUE" *) wire n10883_o;
  (* KEEP="TRUE" *) wire n10884_o;
  (* KEEP="TRUE" *) wire n10885_o;
  (* KEEP="TRUE" *) wire n10886_o;
  (* KEEP="TRUE" *) wire n10887_o;
  (* KEEP="TRUE" *) wire n10888_o;
  (* KEEP="TRUE" *) wire n10889_o;
  (* KEEP="TRUE" *) wire n10890_o;
  (* KEEP="TRUE" *) wire n10891_o;
  (* KEEP="TRUE" *) wire n10892_o;
  (* KEEP="TRUE" *) wire n10893_o;
  (* KEEP="TRUE" *) wire n10894_o;
  (* KEEP="TRUE" *) wire n10895_o;
  (* KEEP="TRUE" *) wire n10896_o;
  (* KEEP="TRUE" *) wire n10897_o;
  (* KEEP="TRUE" *) wire n10898_o;
  (* KEEP="TRUE" *) wire n10899_o;
  (* KEEP="TRUE" *) wire n10900_o;
  (* KEEP="TRUE" *) wire n10901_o;
  (* KEEP="TRUE" *) wire n10902_o;
  (* KEEP="TRUE" *) wire n10903_o;
  (* KEEP="TRUE" *) wire n10904_o;
  (* KEEP="TRUE" *) wire n10905_o;
  (* KEEP="TRUE" *) wire n10906_o;
  (* KEEP="TRUE" *) wire n10907_o;
  (* KEEP="TRUE" *) wire n10908_o;
  (* KEEP="TRUE" *) wire n10909_o;
  (* KEEP="TRUE" *) wire n10910_o;
  (* KEEP="TRUE" *) wire n10911_o;
  (* KEEP="TRUE" *) wire n10912_o;
  (* KEEP="TRUE" *) wire n10913_o;
  (* KEEP="TRUE" *) wire n10914_o;
  (* KEEP="TRUE" *) wire n10915_o;
  (* KEEP="TRUE" *) wire n10916_o;
  (* KEEP="TRUE" *) wire n10917_o;
  (* KEEP="TRUE" *) wire n10918_o;
  (* KEEP="TRUE" *) wire n10919_o;
  (* KEEP="TRUE" *) wire n10920_o;
  (* KEEP="TRUE" *) wire n10921_o;
  (* KEEP="TRUE" *) wire n10922_o;
  (* KEEP="TRUE" *) wire n10923_o;
  (* KEEP="TRUE" *) wire n10924_o;
  (* KEEP="TRUE" *) wire n10925_o;
  (* KEEP="TRUE" *) wire n10926_o;
  (* KEEP="TRUE" *) wire n10927_o;
  (* KEEP="TRUE" *) wire n10928_o;
  (* KEEP="TRUE" *) wire n10929_o;
  (* KEEP="TRUE" *) wire n10930_o;
  (* KEEP="TRUE" *) wire n10931_o;
  (* KEEP="TRUE" *) wire n10932_o;
  (* KEEP="TRUE" *) wire n10933_o;
  (* KEEP="TRUE" *) wire n10934_o;
  (* KEEP="TRUE" *) wire n10935_o;
  (* KEEP="TRUE" *) wire n10936_o;
  (* KEEP="TRUE" *) wire n10937_o;
  (* KEEP="TRUE" *) wire n10938_o;
  (* KEEP="TRUE" *) wire n10939_o;
  (* KEEP="TRUE" *) wire n10940_o;
  (* KEEP="TRUE" *) wire n10941_o;
  (* KEEP="TRUE" *) wire n10942_o;
  (* KEEP="TRUE" *) wire n10943_o;
  (* KEEP="TRUE" *) wire n10944_o;
  (* KEEP="TRUE" *) wire n10945_o;
  (* KEEP="TRUE" *) wire n10946_o;
  (* KEEP="TRUE" *) wire n10947_o;
  (* KEEP="TRUE" *) wire n10948_o;
  (* KEEP="TRUE" *) wire n10949_o;
  (* KEEP="TRUE" *) wire n10950_o;
  (* KEEP="TRUE" *) wire n10951_o;
  (* KEEP="TRUE" *) wire n10952_o;
  (* KEEP="TRUE" *) wire n10953_o;
  (* KEEP="TRUE" *) wire n10954_o;
  (* KEEP="TRUE" *) wire n10955_o;
  (* KEEP="TRUE" *) wire n10956_o;
  (* KEEP="TRUE" *) wire n10957_o;
  (* KEEP="TRUE" *) wire n10958_o;
  (* KEEP="TRUE" *) wire n10959_o;
  (* KEEP="TRUE" *) wire n10960_o;
  (* KEEP="TRUE" *) wire n10961_o;
  (* KEEP="TRUE" *) wire n10962_o;
  (* KEEP="TRUE" *) wire n10963_o;
  (* KEEP="TRUE" *) wire n10964_o;
  (* KEEP="TRUE" *) wire n10965_o;
  (* KEEP="TRUE" *) wire n10966_o;
  (* KEEP="TRUE" *) wire n10967_o;
  (* KEEP="TRUE" *) wire n10968_o;
  (* KEEP="TRUE" *) wire n10969_o;
  (* KEEP="TRUE" *) wire n10970_o;
  (* KEEP="TRUE" *) wire n10971_o;
  (* KEEP="TRUE" *) wire n10972_o;
  (* KEEP="TRUE" *) wire n10973_o;
  (* KEEP="TRUE" *) wire n10974_o;
  (* KEEP="TRUE" *) wire n10975_o;
  (* KEEP="TRUE" *) wire n10976_o;
  (* KEEP="TRUE" *) wire n10977_o;
  (* KEEP="TRUE" *) wire n10978_o;
  (* KEEP="TRUE" *) wire n10979_o;
  (* KEEP="TRUE" *) wire n10980_o;
  (* KEEP="TRUE" *) wire n10981_o;
  (* KEEP="TRUE" *) wire n10982_o;
  (* KEEP="TRUE" *) wire n10983_o;
  (* KEEP="TRUE" *) wire n10984_o;
  (* KEEP="TRUE" *) wire n10985_o;
  (* KEEP="TRUE" *) wire n10986_o;
  (* KEEP="TRUE" *) wire n10987_o;
  (* KEEP="TRUE" *) wire n10988_o;
  (* KEEP="TRUE" *) wire n10989_o;
  (* KEEP="TRUE" *) wire n10990_o;
  (* KEEP="TRUE" *) wire n10991_o;
  (* KEEP="TRUE" *) wire n10992_o;
  (* KEEP="TRUE" *) wire n10993_o;
  (* KEEP="TRUE" *) wire n10994_o;
  (* KEEP="TRUE" *) wire n10995_o;
  (* KEEP="TRUE" *) wire n10996_o;
  (* KEEP="TRUE" *) wire n10997_o;
  (* KEEP="TRUE" *) wire n10998_o;
  (* KEEP="TRUE" *) wire n10999_o;
  (* KEEP="TRUE" *) wire n11000_o;
  (* KEEP="TRUE" *) wire n11001_o;
  (* KEEP="TRUE" *) wire n11002_o;
  (* KEEP="TRUE" *) wire n11003_o;
  (* KEEP="TRUE" *) wire n11004_o;
  (* KEEP="TRUE" *) wire n11005_o;
  (* KEEP="TRUE" *) wire n11006_o;
  (* KEEP="TRUE" *) wire n11007_o;
  (* KEEP="TRUE" *) wire n11008_o;
  (* KEEP="TRUE" *) wire n11009_o;
  (* KEEP="TRUE" *) wire n11010_o;
  (* KEEP="TRUE" *) wire n11011_o;
  (* KEEP="TRUE" *) wire n11012_o;
  (* KEEP="TRUE" *) wire n11013_o;
  (* KEEP="TRUE" *) wire n11014_o;
  (* KEEP="TRUE" *) wire n11015_o;
  (* KEEP="TRUE" *) wire n11016_o;
  (* KEEP="TRUE" *) wire n11017_o;
  (* KEEP="TRUE" *) wire n11018_o;
  (* KEEP="TRUE" *) wire n11019_o;
  (* KEEP="TRUE" *) wire n11020_o;
  (* KEEP="TRUE" *) wire n11021_o;
  (* KEEP="TRUE" *) reg n11022_q;
  assign \output  = n11022_q;
  /* RTL_PUF/vhdl/ro_array.vhd:32:8  */
  assign sortie_ro = n10765_o; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4873_o = enable[0];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n1_ringoscillator_n4874 = inverseur_n1_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n1_ringoscillator (
    .enable(n4873_o),
    .ro_out(inverseur_n1_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4877_o = enable[1];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n2_ringoscillator_n4878 = inverseur_n2_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n2_ringoscillator (
    .enable(n4877_o),
    .ro_out(inverseur_n2_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4881_o = enable[2];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n3_ringoscillator_n4882 = inverseur_n3_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n3_ringoscillator (
    .enable(n4881_o),
    .ro_out(inverseur_n3_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4885_o = enable[3];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n4_ringoscillator_n4886 = inverseur_n4_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n4_ringoscillator (
    .enable(n4885_o),
    .ro_out(inverseur_n4_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4889_o = enable[4];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n5_ringoscillator_n4890 = inverseur_n5_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n5_ringoscillator (
    .enable(n4889_o),
    .ro_out(inverseur_n5_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4893_o = enable[5];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n6_ringoscillator_n4894 = inverseur_n6_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n6_ringoscillator (
    .enable(n4893_o),
    .ro_out(inverseur_n6_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4897_o = enable[6];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n7_ringoscillator_n4898 = inverseur_n7_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n7_ringoscillator (
    .enable(n4897_o),
    .ro_out(inverseur_n7_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4901_o = enable[7];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n8_ringoscillator_n4902 = inverseur_n8_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n8_ringoscillator (
    .enable(n4901_o),
    .ro_out(inverseur_n8_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4905_o = enable[8];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n9_ringoscillator_n4906 = inverseur_n9_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n9_ringoscillator (
    .enable(n4905_o),
    .ro_out(inverseur_n9_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4909_o = enable[9];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n10_ringoscillator_n4910 = inverseur_n10_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n10_ringoscillator (
    .enable(n4909_o),
    .ro_out(inverseur_n10_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4913_o = enable[10];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n11_ringoscillator_n4914 = inverseur_n11_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n11_ringoscillator (
    .enable(n4913_o),
    .ro_out(inverseur_n11_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4917_o = enable[11];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n12_ringoscillator_n4918 = inverseur_n12_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n12_ringoscillator (
    .enable(n4917_o),
    .ro_out(inverseur_n12_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4921_o = enable[12];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n13_ringoscillator_n4922 = inverseur_n13_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n13_ringoscillator (
    .enable(n4921_o),
    .ro_out(inverseur_n13_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4925_o = enable[13];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n14_ringoscillator_n4926 = inverseur_n14_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n14_ringoscillator (
    .enable(n4925_o),
    .ro_out(inverseur_n14_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4929_o = enable[14];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n15_ringoscillator_n4930 = inverseur_n15_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n15_ringoscillator (
    .enable(n4929_o),
    .ro_out(inverseur_n15_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4933_o = enable[15];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n16_ringoscillator_n4934 = inverseur_n16_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n16_ringoscillator (
    .enable(n4933_o),
    .ro_out(inverseur_n16_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4937_o = enable[16];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n17_ringoscillator_n4938 = inverseur_n17_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n17_ringoscillator (
    .enable(n4937_o),
    .ro_out(inverseur_n17_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4941_o = enable[17];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n18_ringoscillator_n4942 = inverseur_n18_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n18_ringoscillator (
    .enable(n4941_o),
    .ro_out(inverseur_n18_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4945_o = enable[18];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n19_ringoscillator_n4946 = inverseur_n19_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n19_ringoscillator (
    .enable(n4945_o),
    .ro_out(inverseur_n19_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4949_o = enable[19];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n20_ringoscillator_n4950 = inverseur_n20_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n20_ringoscillator (
    .enable(n4949_o),
    .ro_out(inverseur_n20_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4953_o = enable[20];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n21_ringoscillator_n4954 = inverseur_n21_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n21_ringoscillator (
    .enable(n4953_o),
    .ro_out(inverseur_n21_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4957_o = enable[21];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n22_ringoscillator_n4958 = inverseur_n22_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n22_ringoscillator (
    .enable(n4957_o),
    .ro_out(inverseur_n22_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4961_o = enable[22];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n23_ringoscillator_n4962 = inverseur_n23_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n23_ringoscillator (
    .enable(n4961_o),
    .ro_out(inverseur_n23_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4965_o = enable[23];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n24_ringoscillator_n4966 = inverseur_n24_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n24_ringoscillator (
    .enable(n4965_o),
    .ro_out(inverseur_n24_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4969_o = enable[24];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n25_ringoscillator_n4970 = inverseur_n25_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n25_ringoscillator (
    .enable(n4969_o),
    .ro_out(inverseur_n25_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4973_o = enable[25];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n26_ringoscillator_n4974 = inverseur_n26_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n26_ringoscillator (
    .enable(n4973_o),
    .ro_out(inverseur_n26_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4977_o = enable[26];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n27_ringoscillator_n4978 = inverseur_n27_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n27_ringoscillator (
    .enable(n4977_o),
    .ro_out(inverseur_n27_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4981_o = enable[27];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n28_ringoscillator_n4982 = inverseur_n28_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n28_ringoscillator (
    .enable(n4981_o),
    .ro_out(inverseur_n28_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4985_o = enable[28];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n29_ringoscillator_n4986 = inverseur_n29_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n29_ringoscillator (
    .enable(n4985_o),
    .ro_out(inverseur_n29_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4989_o = enable[29];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n30_ringoscillator_n4990 = inverseur_n30_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n30_ringoscillator (
    .enable(n4989_o),
    .ro_out(inverseur_n30_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4993_o = enable[30];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n31_ringoscillator_n4994 = inverseur_n31_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n31_ringoscillator (
    .enable(n4993_o),
    .ro_out(inverseur_n31_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n4997_o = enable[31];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n32_ringoscillator_n4998 = inverseur_n32_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n32_ringoscillator (
    .enable(n4997_o),
    .ro_out(inverseur_n32_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5001_o = enable[32];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n33_ringoscillator_n5002 = inverseur_n33_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n33_ringoscillator (
    .enable(n5001_o),
    .ro_out(inverseur_n33_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5005_o = enable[33];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n34_ringoscillator_n5006 = inverseur_n34_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n34_ringoscillator (
    .enable(n5005_o),
    .ro_out(inverseur_n34_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5009_o = enable[34];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n35_ringoscillator_n5010 = inverseur_n35_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n35_ringoscillator (
    .enable(n5009_o),
    .ro_out(inverseur_n35_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5013_o = enable[35];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n36_ringoscillator_n5014 = inverseur_n36_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n36_ringoscillator (
    .enable(n5013_o),
    .ro_out(inverseur_n36_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5017_o = enable[36];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n37_ringoscillator_n5018 = inverseur_n37_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n37_ringoscillator (
    .enable(n5017_o),
    .ro_out(inverseur_n37_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5021_o = enable[37];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n38_ringoscillator_n5022 = inverseur_n38_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n38_ringoscillator (
    .enable(n5021_o),
    .ro_out(inverseur_n38_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5025_o = enable[38];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n39_ringoscillator_n5026 = inverseur_n39_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n39_ringoscillator (
    .enable(n5025_o),
    .ro_out(inverseur_n39_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5029_o = enable[39];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n40_ringoscillator_n5030 = inverseur_n40_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n40_ringoscillator (
    .enable(n5029_o),
    .ro_out(inverseur_n40_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5033_o = enable[40];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n41_ringoscillator_n5034 = inverseur_n41_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n41_ringoscillator (
    .enable(n5033_o),
    .ro_out(inverseur_n41_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5037_o = enable[41];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n42_ringoscillator_n5038 = inverseur_n42_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n42_ringoscillator (
    .enable(n5037_o),
    .ro_out(inverseur_n42_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5041_o = enable[42];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n43_ringoscillator_n5042 = inverseur_n43_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n43_ringoscillator (
    .enable(n5041_o),
    .ro_out(inverseur_n43_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5045_o = enable[43];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n44_ringoscillator_n5046 = inverseur_n44_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n44_ringoscillator (
    .enable(n5045_o),
    .ro_out(inverseur_n44_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5049_o = enable[44];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n45_ringoscillator_n5050 = inverseur_n45_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n45_ringoscillator (
    .enable(n5049_o),
    .ro_out(inverseur_n45_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5053_o = enable[45];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n46_ringoscillator_n5054 = inverseur_n46_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n46_ringoscillator (
    .enable(n5053_o),
    .ro_out(inverseur_n46_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5057_o = enable[46];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n47_ringoscillator_n5058 = inverseur_n47_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n47_ringoscillator (
    .enable(n5057_o),
    .ro_out(inverseur_n47_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5061_o = enable[47];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n48_ringoscillator_n5062 = inverseur_n48_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n48_ringoscillator (
    .enable(n5061_o),
    .ro_out(inverseur_n48_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5065_o = enable[48];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n49_ringoscillator_n5066 = inverseur_n49_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n49_ringoscillator (
    .enable(n5065_o),
    .ro_out(inverseur_n49_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5069_o = enable[49];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n50_ringoscillator_n5070 = inverseur_n50_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n50_ringoscillator (
    .enable(n5069_o),
    .ro_out(inverseur_n50_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5073_o = enable[50];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n51_ringoscillator_n5074 = inverseur_n51_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n51_ringoscillator (
    .enable(n5073_o),
    .ro_out(inverseur_n51_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5077_o = enable[51];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n52_ringoscillator_n5078 = inverseur_n52_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n52_ringoscillator (
    .enable(n5077_o),
    .ro_out(inverseur_n52_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5081_o = enable[52];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n53_ringoscillator_n5082 = inverseur_n53_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n53_ringoscillator (
    .enable(n5081_o),
    .ro_out(inverseur_n53_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5085_o = enable[53];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n54_ringoscillator_n5086 = inverseur_n54_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n54_ringoscillator (
    .enable(n5085_o),
    .ro_out(inverseur_n54_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5089_o = enable[54];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n55_ringoscillator_n5090 = inverseur_n55_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n55_ringoscillator (
    .enable(n5089_o),
    .ro_out(inverseur_n55_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5093_o = enable[55];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n56_ringoscillator_n5094 = inverseur_n56_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n56_ringoscillator (
    .enable(n5093_o),
    .ro_out(inverseur_n56_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5097_o = enable[56];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n57_ringoscillator_n5098 = inverseur_n57_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n57_ringoscillator (
    .enable(n5097_o),
    .ro_out(inverseur_n57_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5101_o = enable[57];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n58_ringoscillator_n5102 = inverseur_n58_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n58_ringoscillator (
    .enable(n5101_o),
    .ro_out(inverseur_n58_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5105_o = enable[58];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n59_ringoscillator_n5106 = inverseur_n59_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n59_ringoscillator (
    .enable(n5105_o),
    .ro_out(inverseur_n59_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5109_o = enable[59];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n60_ringoscillator_n5110 = inverseur_n60_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n60_ringoscillator (
    .enable(n5109_o),
    .ro_out(inverseur_n60_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5113_o = enable[60];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n61_ringoscillator_n5114 = inverseur_n61_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n61_ringoscillator (
    .enable(n5113_o),
    .ro_out(inverseur_n61_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5117_o = enable[61];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n62_ringoscillator_n5118 = inverseur_n62_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n62_ringoscillator (
    .enable(n5117_o),
    .ro_out(inverseur_n62_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5121_o = enable[62];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n63_ringoscillator_n5122 = inverseur_n63_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n63_ringoscillator (
    .enable(n5121_o),
    .ro_out(inverseur_n63_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5125_o = enable[63];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n64_ringoscillator_n5126 = inverseur_n64_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n64_ringoscillator (
    .enable(n5125_o),
    .ro_out(inverseur_n64_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5129_o = enable[64];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n65_ringoscillator_n5130 = inverseur_n65_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n65_ringoscillator (
    .enable(n5129_o),
    .ro_out(inverseur_n65_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5133_o = enable[65];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n66_ringoscillator_n5134 = inverseur_n66_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n66_ringoscillator (
    .enable(n5133_o),
    .ro_out(inverseur_n66_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5137_o = enable[66];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n67_ringoscillator_n5138 = inverseur_n67_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n67_ringoscillator (
    .enable(n5137_o),
    .ro_out(inverseur_n67_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5141_o = enable[67];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n68_ringoscillator_n5142 = inverseur_n68_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n68_ringoscillator (
    .enable(n5141_o),
    .ro_out(inverseur_n68_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5145_o = enable[68];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n69_ringoscillator_n5146 = inverseur_n69_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n69_ringoscillator (
    .enable(n5145_o),
    .ro_out(inverseur_n69_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5149_o = enable[69];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n70_ringoscillator_n5150 = inverseur_n70_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n70_ringoscillator (
    .enable(n5149_o),
    .ro_out(inverseur_n70_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5153_o = enable[70];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n71_ringoscillator_n5154 = inverseur_n71_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n71_ringoscillator (
    .enable(n5153_o),
    .ro_out(inverseur_n71_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5157_o = enable[71];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n72_ringoscillator_n5158 = inverseur_n72_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n72_ringoscillator (
    .enable(n5157_o),
    .ro_out(inverseur_n72_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5161_o = enable[72];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n73_ringoscillator_n5162 = inverseur_n73_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n73_ringoscillator (
    .enable(n5161_o),
    .ro_out(inverseur_n73_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5165_o = enable[73];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n74_ringoscillator_n5166 = inverseur_n74_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n74_ringoscillator (
    .enable(n5165_o),
    .ro_out(inverseur_n74_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5169_o = enable[74];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n75_ringoscillator_n5170 = inverseur_n75_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n75_ringoscillator (
    .enable(n5169_o),
    .ro_out(inverseur_n75_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5173_o = enable[75];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n76_ringoscillator_n5174 = inverseur_n76_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n76_ringoscillator (
    .enable(n5173_o),
    .ro_out(inverseur_n76_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5177_o = enable[76];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n77_ringoscillator_n5178 = inverseur_n77_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n77_ringoscillator (
    .enable(n5177_o),
    .ro_out(inverseur_n77_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5181_o = enable[77];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n78_ringoscillator_n5182 = inverseur_n78_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n78_ringoscillator (
    .enable(n5181_o),
    .ro_out(inverseur_n78_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5185_o = enable[78];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n79_ringoscillator_n5186 = inverseur_n79_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n79_ringoscillator (
    .enable(n5185_o),
    .ro_out(inverseur_n79_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5189_o = enable[79];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n80_ringoscillator_n5190 = inverseur_n80_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n80_ringoscillator (
    .enable(n5189_o),
    .ro_out(inverseur_n80_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5193_o = enable[80];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n81_ringoscillator_n5194 = inverseur_n81_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n81_ringoscillator (
    .enable(n5193_o),
    .ro_out(inverseur_n81_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5197_o = enable[81];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n82_ringoscillator_n5198 = inverseur_n82_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n82_ringoscillator (
    .enable(n5197_o),
    .ro_out(inverseur_n82_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5201_o = enable[82];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n83_ringoscillator_n5202 = inverseur_n83_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n83_ringoscillator (
    .enable(n5201_o),
    .ro_out(inverseur_n83_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5205_o = enable[83];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n84_ringoscillator_n5206 = inverseur_n84_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n84_ringoscillator (
    .enable(n5205_o),
    .ro_out(inverseur_n84_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5209_o = enable[84];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n85_ringoscillator_n5210 = inverseur_n85_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n85_ringoscillator (
    .enable(n5209_o),
    .ro_out(inverseur_n85_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5213_o = enable[85];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n86_ringoscillator_n5214 = inverseur_n86_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n86_ringoscillator (
    .enable(n5213_o),
    .ro_out(inverseur_n86_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5217_o = enable[86];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n87_ringoscillator_n5218 = inverseur_n87_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n87_ringoscillator (
    .enable(n5217_o),
    .ro_out(inverseur_n87_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5221_o = enable[87];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n88_ringoscillator_n5222 = inverseur_n88_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n88_ringoscillator (
    .enable(n5221_o),
    .ro_out(inverseur_n88_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5225_o = enable[88];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n89_ringoscillator_n5226 = inverseur_n89_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n89_ringoscillator (
    .enable(n5225_o),
    .ro_out(inverseur_n89_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5229_o = enable[89];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n90_ringoscillator_n5230 = inverseur_n90_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n90_ringoscillator (
    .enable(n5229_o),
    .ro_out(inverseur_n90_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5233_o = enable[90];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n91_ringoscillator_n5234 = inverseur_n91_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n91_ringoscillator (
    .enable(n5233_o),
    .ro_out(inverseur_n91_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5237_o = enable[91];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n92_ringoscillator_n5238 = inverseur_n92_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n92_ringoscillator (
    .enable(n5237_o),
    .ro_out(inverseur_n92_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5241_o = enable[92];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n93_ringoscillator_n5242 = inverseur_n93_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n93_ringoscillator (
    .enable(n5241_o),
    .ro_out(inverseur_n93_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5245_o = enable[93];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n94_ringoscillator_n5246 = inverseur_n94_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n94_ringoscillator (
    .enable(n5245_o),
    .ro_out(inverseur_n94_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5249_o = enable[94];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n95_ringoscillator_n5250 = inverseur_n95_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n95_ringoscillator (
    .enable(n5249_o),
    .ro_out(inverseur_n95_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5253_o = enable[95];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n96_ringoscillator_n5254 = inverseur_n96_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n96_ringoscillator (
    .enable(n5253_o),
    .ro_out(inverseur_n96_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5257_o = enable[96];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n97_ringoscillator_n5258 = inverseur_n97_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n97_ringoscillator (
    .enable(n5257_o),
    .ro_out(inverseur_n97_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5261_o = enable[97];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n98_ringoscillator_n5262 = inverseur_n98_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n98_ringoscillator (
    .enable(n5261_o),
    .ro_out(inverseur_n98_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5265_o = enable[98];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n99_ringoscillator_n5266 = inverseur_n99_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n99_ringoscillator (
    .enable(n5265_o),
    .ro_out(inverseur_n99_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5269_o = enable[99];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n100_ringoscillator_n5270 = inverseur_n100_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n100_ringoscillator (
    .enable(n5269_o),
    .ro_out(inverseur_n100_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5273_o = enable[100];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n101_ringoscillator_n5274 = inverseur_n101_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n101_ringoscillator (
    .enable(n5273_o),
    .ro_out(inverseur_n101_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5277_o = enable[101];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n102_ringoscillator_n5278 = inverseur_n102_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n102_ringoscillator (
    .enable(n5277_o),
    .ro_out(inverseur_n102_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5281_o = enable[102];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n103_ringoscillator_n5282 = inverseur_n103_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n103_ringoscillator (
    .enable(n5281_o),
    .ro_out(inverseur_n103_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5285_o = enable[103];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n104_ringoscillator_n5286 = inverseur_n104_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n104_ringoscillator (
    .enable(n5285_o),
    .ro_out(inverseur_n104_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5289_o = enable[104];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n105_ringoscillator_n5290 = inverseur_n105_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n105_ringoscillator (
    .enable(n5289_o),
    .ro_out(inverseur_n105_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5293_o = enable[105];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n106_ringoscillator_n5294 = inverseur_n106_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n106_ringoscillator (
    .enable(n5293_o),
    .ro_out(inverseur_n106_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5297_o = enable[106];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n107_ringoscillator_n5298 = inverseur_n107_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n107_ringoscillator (
    .enable(n5297_o),
    .ro_out(inverseur_n107_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5301_o = enable[107];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n108_ringoscillator_n5302 = inverseur_n108_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n108_ringoscillator (
    .enable(n5301_o),
    .ro_out(inverseur_n108_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5305_o = enable[108];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n109_ringoscillator_n5306 = inverseur_n109_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n109_ringoscillator (
    .enable(n5305_o),
    .ro_out(inverseur_n109_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5309_o = enable[109];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n110_ringoscillator_n5310 = inverseur_n110_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n110_ringoscillator (
    .enable(n5309_o),
    .ro_out(inverseur_n110_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5313_o = enable[110];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n111_ringoscillator_n5314 = inverseur_n111_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n111_ringoscillator (
    .enable(n5313_o),
    .ro_out(inverseur_n111_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5317_o = enable[111];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n112_ringoscillator_n5318 = inverseur_n112_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n112_ringoscillator (
    .enable(n5317_o),
    .ro_out(inverseur_n112_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5321_o = enable[112];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n113_ringoscillator_n5322 = inverseur_n113_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n113_ringoscillator (
    .enable(n5321_o),
    .ro_out(inverseur_n113_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5325_o = enable[113];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n114_ringoscillator_n5326 = inverseur_n114_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n114_ringoscillator (
    .enable(n5325_o),
    .ro_out(inverseur_n114_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5329_o = enable[114];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n115_ringoscillator_n5330 = inverseur_n115_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n115_ringoscillator (
    .enable(n5329_o),
    .ro_out(inverseur_n115_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5333_o = enable[115];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n116_ringoscillator_n5334 = inverseur_n116_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n116_ringoscillator (
    .enable(n5333_o),
    .ro_out(inverseur_n116_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5337_o = enable[116];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n117_ringoscillator_n5338 = inverseur_n117_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n117_ringoscillator (
    .enable(n5337_o),
    .ro_out(inverseur_n117_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5341_o = enable[117];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n118_ringoscillator_n5342 = inverseur_n118_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n118_ringoscillator (
    .enable(n5341_o),
    .ro_out(inverseur_n118_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5345_o = enable[118];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n119_ringoscillator_n5346 = inverseur_n119_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n119_ringoscillator (
    .enable(n5345_o),
    .ro_out(inverseur_n119_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5349_o = enable[119];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n120_ringoscillator_n5350 = inverseur_n120_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n120_ringoscillator (
    .enable(n5349_o),
    .ro_out(inverseur_n120_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5353_o = enable[120];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n121_ringoscillator_n5354 = inverseur_n121_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n121_ringoscillator (
    .enable(n5353_o),
    .ro_out(inverseur_n121_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5357_o = enable[121];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n122_ringoscillator_n5358 = inverseur_n122_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n122_ringoscillator (
    .enable(n5357_o),
    .ro_out(inverseur_n122_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5361_o = enable[122];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n123_ringoscillator_n5362 = inverseur_n123_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n123_ringoscillator (
    .enable(n5361_o),
    .ro_out(inverseur_n123_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5365_o = enable[123];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n124_ringoscillator_n5366 = inverseur_n124_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n124_ringoscillator (
    .enable(n5365_o),
    .ro_out(inverseur_n124_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5369_o = enable[124];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n125_ringoscillator_n5370 = inverseur_n125_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n125_ringoscillator (
    .enable(n5369_o),
    .ro_out(inverseur_n125_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5373_o = enable[125];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n126_ringoscillator_n5374 = inverseur_n126_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n126_ringoscillator (
    .enable(n5373_o),
    .ro_out(inverseur_n126_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5377_o = enable[126];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n127_ringoscillator_n5378 = inverseur_n127_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n127_ringoscillator (
    .enable(n5377_o),
    .ro_out(inverseur_n127_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5381_o = enable[127];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n128_ringoscillator_n5382 = inverseur_n128_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n128_ringoscillator (
    .enable(n5381_o),
    .ro_out(inverseur_n128_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5385_o = enable[128];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n129_ringoscillator_n5386 = inverseur_n129_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n129_ringoscillator (
    .enable(n5385_o),
    .ro_out(inverseur_n129_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5389_o = enable[129];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n130_ringoscillator_n5390 = inverseur_n130_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n130_ringoscillator (
    .enable(n5389_o),
    .ro_out(inverseur_n130_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5393_o = enable[130];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n131_ringoscillator_n5394 = inverseur_n131_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n131_ringoscillator (
    .enable(n5393_o),
    .ro_out(inverseur_n131_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5397_o = enable[131];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n132_ringoscillator_n5398 = inverseur_n132_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n132_ringoscillator (
    .enable(n5397_o),
    .ro_out(inverseur_n132_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5401_o = enable[132];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n133_ringoscillator_n5402 = inverseur_n133_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n133_ringoscillator (
    .enable(n5401_o),
    .ro_out(inverseur_n133_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5405_o = enable[133];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n134_ringoscillator_n5406 = inverseur_n134_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n134_ringoscillator (
    .enable(n5405_o),
    .ro_out(inverseur_n134_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5409_o = enable[134];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n135_ringoscillator_n5410 = inverseur_n135_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n135_ringoscillator (
    .enable(n5409_o),
    .ro_out(inverseur_n135_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5413_o = enable[135];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n136_ringoscillator_n5414 = inverseur_n136_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n136_ringoscillator (
    .enable(n5413_o),
    .ro_out(inverseur_n136_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5417_o = enable[136];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n137_ringoscillator_n5418 = inverseur_n137_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n137_ringoscillator (
    .enable(n5417_o),
    .ro_out(inverseur_n137_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5421_o = enable[137];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n138_ringoscillator_n5422 = inverseur_n138_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n138_ringoscillator (
    .enable(n5421_o),
    .ro_out(inverseur_n138_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5425_o = enable[138];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n139_ringoscillator_n5426 = inverseur_n139_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n139_ringoscillator (
    .enable(n5425_o),
    .ro_out(inverseur_n139_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5429_o = enable[139];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n140_ringoscillator_n5430 = inverseur_n140_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n140_ringoscillator (
    .enable(n5429_o),
    .ro_out(inverseur_n140_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5433_o = enable[140];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n141_ringoscillator_n5434 = inverseur_n141_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n141_ringoscillator (
    .enable(n5433_o),
    .ro_out(inverseur_n141_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5437_o = enable[141];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n142_ringoscillator_n5438 = inverseur_n142_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n142_ringoscillator (
    .enable(n5437_o),
    .ro_out(inverseur_n142_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5441_o = enable[142];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n143_ringoscillator_n5442 = inverseur_n143_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n143_ringoscillator (
    .enable(n5441_o),
    .ro_out(inverseur_n143_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5445_o = enable[143];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n144_ringoscillator_n5446 = inverseur_n144_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n144_ringoscillator (
    .enable(n5445_o),
    .ro_out(inverseur_n144_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5449_o = enable[144];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n145_ringoscillator_n5450 = inverseur_n145_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n145_ringoscillator (
    .enable(n5449_o),
    .ro_out(inverseur_n145_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5453_o = enable[145];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n146_ringoscillator_n5454 = inverseur_n146_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n146_ringoscillator (
    .enable(n5453_o),
    .ro_out(inverseur_n146_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5457_o = enable[146];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n147_ringoscillator_n5458 = inverseur_n147_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n147_ringoscillator (
    .enable(n5457_o),
    .ro_out(inverseur_n147_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5461_o = enable[147];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n148_ringoscillator_n5462 = inverseur_n148_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n148_ringoscillator (
    .enable(n5461_o),
    .ro_out(inverseur_n148_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5465_o = enable[148];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n149_ringoscillator_n5466 = inverseur_n149_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n149_ringoscillator (
    .enable(n5465_o),
    .ro_out(inverseur_n149_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5469_o = enable[149];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n150_ringoscillator_n5470 = inverseur_n150_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n150_ringoscillator (
    .enable(n5469_o),
    .ro_out(inverseur_n150_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5473_o = enable[150];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n151_ringoscillator_n5474 = inverseur_n151_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n151_ringoscillator (
    .enable(n5473_o),
    .ro_out(inverseur_n151_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5477_o = enable[151];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n152_ringoscillator_n5478 = inverseur_n152_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n152_ringoscillator (
    .enable(n5477_o),
    .ro_out(inverseur_n152_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5481_o = enable[152];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n153_ringoscillator_n5482 = inverseur_n153_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n153_ringoscillator (
    .enable(n5481_o),
    .ro_out(inverseur_n153_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5485_o = enable[153];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n154_ringoscillator_n5486 = inverseur_n154_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n154_ringoscillator (
    .enable(n5485_o),
    .ro_out(inverseur_n154_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5489_o = enable[154];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n155_ringoscillator_n5490 = inverseur_n155_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n155_ringoscillator (
    .enable(n5489_o),
    .ro_out(inverseur_n155_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5493_o = enable[155];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n156_ringoscillator_n5494 = inverseur_n156_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n156_ringoscillator (
    .enable(n5493_o),
    .ro_out(inverseur_n156_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5497_o = enable[156];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n157_ringoscillator_n5498 = inverseur_n157_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n157_ringoscillator (
    .enable(n5497_o),
    .ro_out(inverseur_n157_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5501_o = enable[157];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n158_ringoscillator_n5502 = inverseur_n158_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n158_ringoscillator (
    .enable(n5501_o),
    .ro_out(inverseur_n158_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5505_o = enable[158];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n159_ringoscillator_n5506 = inverseur_n159_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n159_ringoscillator (
    .enable(n5505_o),
    .ro_out(inverseur_n159_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5509_o = enable[159];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n160_ringoscillator_n5510 = inverseur_n160_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n160_ringoscillator (
    .enable(n5509_o),
    .ro_out(inverseur_n160_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5513_o = enable[160];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n161_ringoscillator_n5514 = inverseur_n161_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n161_ringoscillator (
    .enable(n5513_o),
    .ro_out(inverseur_n161_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5517_o = enable[161];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n162_ringoscillator_n5518 = inverseur_n162_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n162_ringoscillator (
    .enable(n5517_o),
    .ro_out(inverseur_n162_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5521_o = enable[162];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n163_ringoscillator_n5522 = inverseur_n163_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n163_ringoscillator (
    .enable(n5521_o),
    .ro_out(inverseur_n163_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5525_o = enable[163];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n164_ringoscillator_n5526 = inverseur_n164_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n164_ringoscillator (
    .enable(n5525_o),
    .ro_out(inverseur_n164_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5529_o = enable[164];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n165_ringoscillator_n5530 = inverseur_n165_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n165_ringoscillator (
    .enable(n5529_o),
    .ro_out(inverseur_n165_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5533_o = enable[165];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n166_ringoscillator_n5534 = inverseur_n166_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n166_ringoscillator (
    .enable(n5533_o),
    .ro_out(inverseur_n166_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5537_o = enable[166];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n167_ringoscillator_n5538 = inverseur_n167_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n167_ringoscillator (
    .enable(n5537_o),
    .ro_out(inverseur_n167_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5541_o = enable[167];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n168_ringoscillator_n5542 = inverseur_n168_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n168_ringoscillator (
    .enable(n5541_o),
    .ro_out(inverseur_n168_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5545_o = enable[168];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n169_ringoscillator_n5546 = inverseur_n169_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n169_ringoscillator (
    .enable(n5545_o),
    .ro_out(inverseur_n169_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5549_o = enable[169];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n170_ringoscillator_n5550 = inverseur_n170_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n170_ringoscillator (
    .enable(n5549_o),
    .ro_out(inverseur_n170_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5553_o = enable[170];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n171_ringoscillator_n5554 = inverseur_n171_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n171_ringoscillator (
    .enable(n5553_o),
    .ro_out(inverseur_n171_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5557_o = enable[171];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n172_ringoscillator_n5558 = inverseur_n172_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n172_ringoscillator (
    .enable(n5557_o),
    .ro_out(inverseur_n172_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5561_o = enable[172];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n173_ringoscillator_n5562 = inverseur_n173_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n173_ringoscillator (
    .enable(n5561_o),
    .ro_out(inverseur_n173_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5565_o = enable[173];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n174_ringoscillator_n5566 = inverseur_n174_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n174_ringoscillator (
    .enable(n5565_o),
    .ro_out(inverseur_n174_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5569_o = enable[174];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n175_ringoscillator_n5570 = inverseur_n175_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n175_ringoscillator (
    .enable(n5569_o),
    .ro_out(inverseur_n175_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5573_o = enable[175];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n176_ringoscillator_n5574 = inverseur_n176_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n176_ringoscillator (
    .enable(n5573_o),
    .ro_out(inverseur_n176_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5577_o = enable[176];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n177_ringoscillator_n5578 = inverseur_n177_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n177_ringoscillator (
    .enable(n5577_o),
    .ro_out(inverseur_n177_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5581_o = enable[177];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n178_ringoscillator_n5582 = inverseur_n178_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n178_ringoscillator (
    .enable(n5581_o),
    .ro_out(inverseur_n178_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5585_o = enable[178];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n179_ringoscillator_n5586 = inverseur_n179_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n179_ringoscillator (
    .enable(n5585_o),
    .ro_out(inverseur_n179_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5589_o = enable[179];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n180_ringoscillator_n5590 = inverseur_n180_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n180_ringoscillator (
    .enable(n5589_o),
    .ro_out(inverseur_n180_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5593_o = enable[180];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n181_ringoscillator_n5594 = inverseur_n181_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n181_ringoscillator (
    .enable(n5593_o),
    .ro_out(inverseur_n181_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5597_o = enable[181];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n182_ringoscillator_n5598 = inverseur_n182_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n182_ringoscillator (
    .enable(n5597_o),
    .ro_out(inverseur_n182_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5601_o = enable[182];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n183_ringoscillator_n5602 = inverseur_n183_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n183_ringoscillator (
    .enable(n5601_o),
    .ro_out(inverseur_n183_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5605_o = enable[183];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n184_ringoscillator_n5606 = inverseur_n184_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n184_ringoscillator (
    .enable(n5605_o),
    .ro_out(inverseur_n184_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5609_o = enable[184];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n185_ringoscillator_n5610 = inverseur_n185_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n185_ringoscillator (
    .enable(n5609_o),
    .ro_out(inverseur_n185_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5613_o = enable[185];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n186_ringoscillator_n5614 = inverseur_n186_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n186_ringoscillator (
    .enable(n5613_o),
    .ro_out(inverseur_n186_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5617_o = enable[186];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n187_ringoscillator_n5618 = inverseur_n187_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n187_ringoscillator (
    .enable(n5617_o),
    .ro_out(inverseur_n187_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5621_o = enable[187];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n188_ringoscillator_n5622 = inverseur_n188_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n188_ringoscillator (
    .enable(n5621_o),
    .ro_out(inverseur_n188_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5625_o = enable[188];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n189_ringoscillator_n5626 = inverseur_n189_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n189_ringoscillator (
    .enable(n5625_o),
    .ro_out(inverseur_n189_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5629_o = enable[189];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n190_ringoscillator_n5630 = inverseur_n190_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n190_ringoscillator (
    .enable(n5629_o),
    .ro_out(inverseur_n190_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5633_o = enable[190];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n191_ringoscillator_n5634 = inverseur_n191_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n191_ringoscillator (
    .enable(n5633_o),
    .ro_out(inverseur_n191_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5637_o = enable[191];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n192_ringoscillator_n5638 = inverseur_n192_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n192_ringoscillator (
    .enable(n5637_o),
    .ro_out(inverseur_n192_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5641_o = enable[192];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n193_ringoscillator_n5642 = inverseur_n193_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n193_ringoscillator (
    .enable(n5641_o),
    .ro_out(inverseur_n193_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5645_o = enable[193];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n194_ringoscillator_n5646 = inverseur_n194_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n194_ringoscillator (
    .enable(n5645_o),
    .ro_out(inverseur_n194_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5649_o = enable[194];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n195_ringoscillator_n5650 = inverseur_n195_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n195_ringoscillator (
    .enable(n5649_o),
    .ro_out(inverseur_n195_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5653_o = enable[195];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n196_ringoscillator_n5654 = inverseur_n196_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n196_ringoscillator (
    .enable(n5653_o),
    .ro_out(inverseur_n196_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5657_o = enable[196];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n197_ringoscillator_n5658 = inverseur_n197_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n197_ringoscillator (
    .enable(n5657_o),
    .ro_out(inverseur_n197_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5661_o = enable[197];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n198_ringoscillator_n5662 = inverseur_n198_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n198_ringoscillator (
    .enable(n5661_o),
    .ro_out(inverseur_n198_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5665_o = enable[198];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n199_ringoscillator_n5666 = inverseur_n199_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n199_ringoscillator (
    .enable(n5665_o),
    .ro_out(inverseur_n199_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5669_o = enable[199];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n200_ringoscillator_n5670 = inverseur_n200_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n200_ringoscillator (
    .enable(n5669_o),
    .ro_out(inverseur_n200_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5673_o = enable[200];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n201_ringoscillator_n5674 = inverseur_n201_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n201_ringoscillator (
    .enable(n5673_o),
    .ro_out(inverseur_n201_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5677_o = enable[201];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n202_ringoscillator_n5678 = inverseur_n202_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n202_ringoscillator (
    .enable(n5677_o),
    .ro_out(inverseur_n202_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5681_o = enable[202];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n203_ringoscillator_n5682 = inverseur_n203_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n203_ringoscillator (
    .enable(n5681_o),
    .ro_out(inverseur_n203_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5685_o = enable[203];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n204_ringoscillator_n5686 = inverseur_n204_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n204_ringoscillator (
    .enable(n5685_o),
    .ro_out(inverseur_n204_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5689_o = enable[204];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n205_ringoscillator_n5690 = inverseur_n205_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n205_ringoscillator (
    .enable(n5689_o),
    .ro_out(inverseur_n205_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5693_o = enable[205];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n206_ringoscillator_n5694 = inverseur_n206_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n206_ringoscillator (
    .enable(n5693_o),
    .ro_out(inverseur_n206_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5697_o = enable[206];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n207_ringoscillator_n5698 = inverseur_n207_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n207_ringoscillator (
    .enable(n5697_o),
    .ro_out(inverseur_n207_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5701_o = enable[207];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n208_ringoscillator_n5702 = inverseur_n208_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n208_ringoscillator (
    .enable(n5701_o),
    .ro_out(inverseur_n208_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5705_o = enable[208];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n209_ringoscillator_n5706 = inverseur_n209_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n209_ringoscillator (
    .enable(n5705_o),
    .ro_out(inverseur_n209_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5709_o = enable[209];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n210_ringoscillator_n5710 = inverseur_n210_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n210_ringoscillator (
    .enable(n5709_o),
    .ro_out(inverseur_n210_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5713_o = enable[210];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n211_ringoscillator_n5714 = inverseur_n211_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n211_ringoscillator (
    .enable(n5713_o),
    .ro_out(inverseur_n211_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5717_o = enable[211];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n212_ringoscillator_n5718 = inverseur_n212_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n212_ringoscillator (
    .enable(n5717_o),
    .ro_out(inverseur_n212_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5721_o = enable[212];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n213_ringoscillator_n5722 = inverseur_n213_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n213_ringoscillator (
    .enable(n5721_o),
    .ro_out(inverseur_n213_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5725_o = enable[213];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n214_ringoscillator_n5726 = inverseur_n214_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n214_ringoscillator (
    .enable(n5725_o),
    .ro_out(inverseur_n214_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5729_o = enable[214];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n215_ringoscillator_n5730 = inverseur_n215_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n215_ringoscillator (
    .enable(n5729_o),
    .ro_out(inverseur_n215_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5733_o = enable[215];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n216_ringoscillator_n5734 = inverseur_n216_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n216_ringoscillator (
    .enable(n5733_o),
    .ro_out(inverseur_n216_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5737_o = enable[216];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n217_ringoscillator_n5738 = inverseur_n217_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n217_ringoscillator (
    .enable(n5737_o),
    .ro_out(inverseur_n217_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5741_o = enable[217];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n218_ringoscillator_n5742 = inverseur_n218_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n218_ringoscillator (
    .enable(n5741_o),
    .ro_out(inverseur_n218_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5745_o = enable[218];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n219_ringoscillator_n5746 = inverseur_n219_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n219_ringoscillator (
    .enable(n5745_o),
    .ro_out(inverseur_n219_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5749_o = enable[219];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n220_ringoscillator_n5750 = inverseur_n220_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n220_ringoscillator (
    .enable(n5749_o),
    .ro_out(inverseur_n220_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5753_o = enable[220];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n221_ringoscillator_n5754 = inverseur_n221_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n221_ringoscillator (
    .enable(n5753_o),
    .ro_out(inverseur_n221_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5757_o = enable[221];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n222_ringoscillator_n5758 = inverseur_n222_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n222_ringoscillator (
    .enable(n5757_o),
    .ro_out(inverseur_n222_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5761_o = enable[222];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n223_ringoscillator_n5762 = inverseur_n223_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n223_ringoscillator (
    .enable(n5761_o),
    .ro_out(inverseur_n223_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5765_o = enable[223];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n224_ringoscillator_n5766 = inverseur_n224_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n224_ringoscillator (
    .enable(n5765_o),
    .ro_out(inverseur_n224_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5769_o = enable[224];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n225_ringoscillator_n5770 = inverseur_n225_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n225_ringoscillator (
    .enable(n5769_o),
    .ro_out(inverseur_n225_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5773_o = enable[225];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n226_ringoscillator_n5774 = inverseur_n226_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n226_ringoscillator (
    .enable(n5773_o),
    .ro_out(inverseur_n226_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5777_o = enable[226];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n227_ringoscillator_n5778 = inverseur_n227_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n227_ringoscillator (
    .enable(n5777_o),
    .ro_out(inverseur_n227_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5781_o = enable[227];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n228_ringoscillator_n5782 = inverseur_n228_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n228_ringoscillator (
    .enable(n5781_o),
    .ro_out(inverseur_n228_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5785_o = enable[228];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n229_ringoscillator_n5786 = inverseur_n229_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n229_ringoscillator (
    .enable(n5785_o),
    .ro_out(inverseur_n229_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5789_o = enable[229];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n230_ringoscillator_n5790 = inverseur_n230_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n230_ringoscillator (
    .enable(n5789_o),
    .ro_out(inverseur_n230_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5793_o = enable[230];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n231_ringoscillator_n5794 = inverseur_n231_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n231_ringoscillator (
    .enable(n5793_o),
    .ro_out(inverseur_n231_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5797_o = enable[231];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n232_ringoscillator_n5798 = inverseur_n232_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n232_ringoscillator (
    .enable(n5797_o),
    .ro_out(inverseur_n232_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5801_o = enable[232];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n233_ringoscillator_n5802 = inverseur_n233_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n233_ringoscillator (
    .enable(n5801_o),
    .ro_out(inverseur_n233_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5805_o = enable[233];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n234_ringoscillator_n5806 = inverseur_n234_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n234_ringoscillator (
    .enable(n5805_o),
    .ro_out(inverseur_n234_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5809_o = enable[234];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n235_ringoscillator_n5810 = inverseur_n235_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n235_ringoscillator (
    .enable(n5809_o),
    .ro_out(inverseur_n235_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5813_o = enable[235];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n236_ringoscillator_n5814 = inverseur_n236_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n236_ringoscillator (
    .enable(n5813_o),
    .ro_out(inverseur_n236_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5817_o = enable[236];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n237_ringoscillator_n5818 = inverseur_n237_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n237_ringoscillator (
    .enable(n5817_o),
    .ro_out(inverseur_n237_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5821_o = enable[237];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n238_ringoscillator_n5822 = inverseur_n238_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n238_ringoscillator (
    .enable(n5821_o),
    .ro_out(inverseur_n238_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5825_o = enable[238];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n239_ringoscillator_n5826 = inverseur_n239_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n239_ringoscillator (
    .enable(n5825_o),
    .ro_out(inverseur_n239_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5829_o = enable[239];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n240_ringoscillator_n5830 = inverseur_n240_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n240_ringoscillator (
    .enable(n5829_o),
    .ro_out(inverseur_n240_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5833_o = enable[240];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n241_ringoscillator_n5834 = inverseur_n241_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n241_ringoscillator (
    .enable(n5833_o),
    .ro_out(inverseur_n241_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5837_o = enable[241];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n242_ringoscillator_n5838 = inverseur_n242_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n242_ringoscillator (
    .enable(n5837_o),
    .ro_out(inverseur_n242_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5841_o = enable[242];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n243_ringoscillator_n5842 = inverseur_n243_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n243_ringoscillator (
    .enable(n5841_o),
    .ro_out(inverseur_n243_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5845_o = enable[243];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n244_ringoscillator_n5846 = inverseur_n244_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n244_ringoscillator (
    .enable(n5845_o),
    .ro_out(inverseur_n244_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5849_o = enable[244];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n245_ringoscillator_n5850 = inverseur_n245_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n245_ringoscillator (
    .enable(n5849_o),
    .ro_out(inverseur_n245_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5853_o = enable[245];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n246_ringoscillator_n5854 = inverseur_n246_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n246_ringoscillator (
    .enable(n5853_o),
    .ro_out(inverseur_n246_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5857_o = enable[246];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n247_ringoscillator_n5858 = inverseur_n247_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n247_ringoscillator (
    .enable(n5857_o),
    .ro_out(inverseur_n247_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5861_o = enable[247];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n248_ringoscillator_n5862 = inverseur_n248_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n248_ringoscillator (
    .enable(n5861_o),
    .ro_out(inverseur_n248_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5865_o = enable[248];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n249_ringoscillator_n5866 = inverseur_n249_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n249_ringoscillator (
    .enable(n5865_o),
    .ro_out(inverseur_n249_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5869_o = enable[249];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n250_ringoscillator_n5870 = inverseur_n250_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n250_ringoscillator (
    .enable(n5869_o),
    .ro_out(inverseur_n250_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5873_o = enable[250];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n251_ringoscillator_n5874 = inverseur_n251_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n251_ringoscillator (
    .enable(n5873_o),
    .ro_out(inverseur_n251_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5877_o = enable[251];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n252_ringoscillator_n5878 = inverseur_n252_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n252_ringoscillator (
    .enable(n5877_o),
    .ro_out(inverseur_n252_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5881_o = enable[252];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n253_ringoscillator_n5882 = inverseur_n253_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n253_ringoscillator (
    .enable(n5881_o),
    .ro_out(inverseur_n253_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5885_o = enable[253];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n254_ringoscillator_n5886 = inverseur_n254_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n254_ringoscillator (
    .enable(n5885_o),
    .ro_out(inverseur_n254_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5889_o = enable[254];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n255_ringoscillator_n5890 = inverseur_n255_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n255_ringoscillator (
    .enable(n5889_o),
    .ro_out(inverseur_n255_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:39:31  */
  assign n5893_o = enable[255];
  /* RTL_PUF/vhdl/ro_array.vhd:40:25  */
  assign inverseur_n256_ringoscillator_n5894 = inverseur_n256_ringoscillator_ro_out; // (signal)
  /* RTL_PUF/vhdl/ro_array.vhd:37:5  */
  ring_oscillator inverseur_n256_ringoscillator (
    .enable(n5893_o),
    .ro_out(inverseur_n256_ringoscillator_ro_out));
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n5902_o = challenge == 8'b00000000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n5903_o = sortie_ro[0];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5913_o = n5902_o ? 1'b0 : 1'b1;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n5916_o = challenge == 8'b00000001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n5917_o = sortie_ro[1];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5918_o = n5929_o ? n5917_o : n5903_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5920_o = n5931_o ? 1'b1 : 1'b1;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5924_o = n5932_o ? 1'b0 : n5913_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5925_o = n5913_o & n5916_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5927_o = n5913_o & n5916_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5928_o = n5913_o & n5916_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5929_o = n5925_o & n5913_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5931_o = n5927_o & n5913_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5932_o = n5928_o & n5913_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n5934_o = challenge == 8'b00000010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n5935_o = sortie_ro[2];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5936_o = n5947_o ? n5935_o : n5918_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5938_o = n5949_o ? 1'b1 : n5920_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5942_o = n5950_o ? 1'b0 : n5924_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5943_o = n5924_o & n5934_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5945_o = n5924_o & n5934_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5946_o = n5924_o & n5934_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5947_o = n5943_o & n5924_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5949_o = n5945_o & n5924_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5950_o = n5946_o & n5924_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n5952_o = challenge == 8'b00000011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n5953_o = sortie_ro[3];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5954_o = n5965_o ? n5953_o : n5936_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5956_o = n5967_o ? 1'b1 : n5938_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5960_o = n5968_o ? 1'b0 : n5942_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5961_o = n5942_o & n5952_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5963_o = n5942_o & n5952_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5964_o = n5942_o & n5952_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5965_o = n5961_o & n5942_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5967_o = n5963_o & n5942_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5968_o = n5964_o & n5942_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n5970_o = challenge == 8'b00000100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n5971_o = sortie_ro[4];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5972_o = n5983_o ? n5971_o : n5954_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5974_o = n5985_o ? 1'b1 : n5956_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5978_o = n5986_o ? 1'b0 : n5960_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5979_o = n5960_o & n5970_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5981_o = n5960_o & n5970_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5982_o = n5960_o & n5970_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5983_o = n5979_o & n5960_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5985_o = n5981_o & n5960_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5986_o = n5982_o & n5960_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n5988_o = challenge == 8'b00000101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n5989_o = sortie_ro[5];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5990_o = n6001_o ? n5989_o : n5972_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5992_o = n6003_o ? 1'b1 : n5974_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5996_o = n6004_o ? 1'b0 : n5978_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5997_o = n5978_o & n5988_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n5999_o = n5978_o & n5988_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6000_o = n5978_o & n5988_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6001_o = n5997_o & n5978_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6003_o = n5999_o & n5978_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6004_o = n6000_o & n5978_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6006_o = challenge == 8'b00000110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6007_o = sortie_ro[6];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6008_o = n6019_o ? n6007_o : n5990_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6010_o = n6021_o ? 1'b1 : n5992_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6014_o = n6022_o ? 1'b0 : n5996_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6015_o = n5996_o & n6006_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6017_o = n5996_o & n6006_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6018_o = n5996_o & n6006_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6019_o = n6015_o & n5996_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6021_o = n6017_o & n5996_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6022_o = n6018_o & n5996_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6024_o = challenge == 8'b00000111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6025_o = sortie_ro[7];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6026_o = n6037_o ? n6025_o : n6008_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6028_o = n6039_o ? 1'b1 : n6010_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6032_o = n6040_o ? 1'b0 : n6014_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6033_o = n6014_o & n6024_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6035_o = n6014_o & n6024_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6036_o = n6014_o & n6024_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6037_o = n6033_o & n6014_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6039_o = n6035_o & n6014_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6040_o = n6036_o & n6014_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6042_o = challenge == 8'b00001000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6043_o = sortie_ro[8];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6044_o = n6055_o ? n6043_o : n6026_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6046_o = n6057_o ? 1'b1 : n6028_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6050_o = n6058_o ? 1'b0 : n6032_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6051_o = n6032_o & n6042_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6053_o = n6032_o & n6042_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6054_o = n6032_o & n6042_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6055_o = n6051_o & n6032_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6057_o = n6053_o & n6032_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6058_o = n6054_o & n6032_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6060_o = challenge == 8'b00001001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6061_o = sortie_ro[9];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6062_o = n6073_o ? n6061_o : n6044_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6064_o = n6075_o ? 1'b1 : n6046_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6068_o = n6076_o ? 1'b0 : n6050_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6069_o = n6050_o & n6060_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6071_o = n6050_o & n6060_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6072_o = n6050_o & n6060_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6073_o = n6069_o & n6050_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6075_o = n6071_o & n6050_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6076_o = n6072_o & n6050_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6078_o = challenge == 8'b00001010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6079_o = sortie_ro[10];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6080_o = n6091_o ? n6079_o : n6062_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6082_o = n6093_o ? 1'b1 : n6064_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6086_o = n6094_o ? 1'b0 : n6068_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6087_o = n6068_o & n6078_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6089_o = n6068_o & n6078_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6090_o = n6068_o & n6078_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6091_o = n6087_o & n6068_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6093_o = n6089_o & n6068_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6094_o = n6090_o & n6068_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6096_o = challenge == 8'b00001011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6097_o = sortie_ro[11];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6098_o = n6109_o ? n6097_o : n6080_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6100_o = n6111_o ? 1'b1 : n6082_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6104_o = n6112_o ? 1'b0 : n6086_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6105_o = n6086_o & n6096_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6107_o = n6086_o & n6096_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6108_o = n6086_o & n6096_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6109_o = n6105_o & n6086_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6111_o = n6107_o & n6086_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6112_o = n6108_o & n6086_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6114_o = challenge == 8'b00001100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6115_o = sortie_ro[12];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6116_o = n6127_o ? n6115_o : n6098_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6118_o = n6129_o ? 1'b1 : n6100_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6122_o = n6130_o ? 1'b0 : n6104_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6123_o = n6104_o & n6114_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6125_o = n6104_o & n6114_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6126_o = n6104_o & n6114_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6127_o = n6123_o & n6104_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6129_o = n6125_o & n6104_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6130_o = n6126_o & n6104_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6132_o = challenge == 8'b00001101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6133_o = sortie_ro[13];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6134_o = n6145_o ? n6133_o : n6116_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6136_o = n6147_o ? 1'b1 : n6118_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6140_o = n6148_o ? 1'b0 : n6122_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6141_o = n6122_o & n6132_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6143_o = n6122_o & n6132_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6144_o = n6122_o & n6132_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6145_o = n6141_o & n6122_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6147_o = n6143_o & n6122_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6148_o = n6144_o & n6122_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6150_o = challenge == 8'b00001110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6151_o = sortie_ro[14];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6152_o = n6163_o ? n6151_o : n6134_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6154_o = n6165_o ? 1'b1 : n6136_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6158_o = n6166_o ? 1'b0 : n6140_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6159_o = n6140_o & n6150_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6161_o = n6140_o & n6150_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6162_o = n6140_o & n6150_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6163_o = n6159_o & n6140_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6165_o = n6161_o & n6140_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6166_o = n6162_o & n6140_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6168_o = challenge == 8'b00001111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6169_o = sortie_ro[15];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6170_o = n6181_o ? n6169_o : n6152_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6172_o = n6183_o ? 1'b1 : n6154_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6176_o = n6184_o ? 1'b0 : n6158_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6177_o = n6158_o & n6168_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6179_o = n6158_o & n6168_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6180_o = n6158_o & n6168_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6181_o = n6177_o & n6158_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6183_o = n6179_o & n6158_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6184_o = n6180_o & n6158_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6186_o = challenge == 8'b00010000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6187_o = sortie_ro[16];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6188_o = n6199_o ? n6187_o : n6170_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6190_o = n6201_o ? 1'b1 : n6172_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6194_o = n6202_o ? 1'b0 : n6176_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6195_o = n6176_o & n6186_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6197_o = n6176_o & n6186_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6198_o = n6176_o & n6186_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6199_o = n6195_o & n6176_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6201_o = n6197_o & n6176_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6202_o = n6198_o & n6176_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6204_o = challenge == 8'b00010001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6205_o = sortie_ro[17];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6206_o = n6217_o ? n6205_o : n6188_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6208_o = n6219_o ? 1'b1 : n6190_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6212_o = n6220_o ? 1'b0 : n6194_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6213_o = n6194_o & n6204_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6215_o = n6194_o & n6204_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6216_o = n6194_o & n6204_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6217_o = n6213_o & n6194_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6219_o = n6215_o & n6194_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6220_o = n6216_o & n6194_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6222_o = challenge == 8'b00010010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6223_o = sortie_ro[18];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6224_o = n6235_o ? n6223_o : n6206_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6226_o = n6237_o ? 1'b1 : n6208_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6230_o = n6238_o ? 1'b0 : n6212_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6231_o = n6212_o & n6222_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6233_o = n6212_o & n6222_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6234_o = n6212_o & n6222_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6235_o = n6231_o & n6212_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6237_o = n6233_o & n6212_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6238_o = n6234_o & n6212_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6240_o = challenge == 8'b00010011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6241_o = sortie_ro[19];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6242_o = n6253_o ? n6241_o : n6224_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6244_o = n6255_o ? 1'b1 : n6226_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6248_o = n6256_o ? 1'b0 : n6230_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6249_o = n6230_o & n6240_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6251_o = n6230_o & n6240_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6252_o = n6230_o & n6240_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6253_o = n6249_o & n6230_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6255_o = n6251_o & n6230_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6256_o = n6252_o & n6230_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6258_o = challenge == 8'b00010100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6259_o = sortie_ro[20];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6260_o = n6271_o ? n6259_o : n6242_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6262_o = n6273_o ? 1'b1 : n6244_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6266_o = n6274_o ? 1'b0 : n6248_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6267_o = n6248_o & n6258_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6269_o = n6248_o & n6258_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6270_o = n6248_o & n6258_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6271_o = n6267_o & n6248_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6273_o = n6269_o & n6248_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6274_o = n6270_o & n6248_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6276_o = challenge == 8'b00010101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6277_o = sortie_ro[21];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6278_o = n6289_o ? n6277_o : n6260_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6280_o = n6291_o ? 1'b1 : n6262_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6284_o = n6292_o ? 1'b0 : n6266_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6285_o = n6266_o & n6276_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6287_o = n6266_o & n6276_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6288_o = n6266_o & n6276_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6289_o = n6285_o & n6266_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6291_o = n6287_o & n6266_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6292_o = n6288_o & n6266_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6294_o = challenge == 8'b00010110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6295_o = sortie_ro[22];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6296_o = n6307_o ? n6295_o : n6278_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6298_o = n6309_o ? 1'b1 : n6280_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6302_o = n6310_o ? 1'b0 : n6284_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6303_o = n6284_o & n6294_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6305_o = n6284_o & n6294_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6306_o = n6284_o & n6294_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6307_o = n6303_o & n6284_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6309_o = n6305_o & n6284_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6310_o = n6306_o & n6284_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6312_o = challenge == 8'b00010111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6313_o = sortie_ro[23];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6314_o = n6325_o ? n6313_o : n6296_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6316_o = n6327_o ? 1'b1 : n6298_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6320_o = n6328_o ? 1'b0 : n6302_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6321_o = n6302_o & n6312_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6323_o = n6302_o & n6312_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6324_o = n6302_o & n6312_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6325_o = n6321_o & n6302_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6327_o = n6323_o & n6302_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6328_o = n6324_o & n6302_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6330_o = challenge == 8'b00011000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6331_o = sortie_ro[24];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6332_o = n6343_o ? n6331_o : n6314_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6334_o = n6345_o ? 1'b1 : n6316_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6338_o = n6346_o ? 1'b0 : n6320_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6339_o = n6320_o & n6330_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6341_o = n6320_o & n6330_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6342_o = n6320_o & n6330_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6343_o = n6339_o & n6320_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6345_o = n6341_o & n6320_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6346_o = n6342_o & n6320_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6348_o = challenge == 8'b00011001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6349_o = sortie_ro[25];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6350_o = n6361_o ? n6349_o : n6332_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6352_o = n6363_o ? 1'b1 : n6334_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6356_o = n6364_o ? 1'b0 : n6338_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6357_o = n6338_o & n6348_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6359_o = n6338_o & n6348_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6360_o = n6338_o & n6348_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6361_o = n6357_o & n6338_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6363_o = n6359_o & n6338_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6364_o = n6360_o & n6338_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6366_o = challenge == 8'b00011010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6367_o = sortie_ro[26];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6368_o = n6379_o ? n6367_o : n6350_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6370_o = n6381_o ? 1'b1 : n6352_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6374_o = n6382_o ? 1'b0 : n6356_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6375_o = n6356_o & n6366_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6377_o = n6356_o & n6366_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6378_o = n6356_o & n6366_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6379_o = n6375_o & n6356_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6381_o = n6377_o & n6356_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6382_o = n6378_o & n6356_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6384_o = challenge == 8'b00011011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6385_o = sortie_ro[27];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6386_o = n6397_o ? n6385_o : n6368_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6388_o = n6399_o ? 1'b1 : n6370_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6392_o = n6400_o ? 1'b0 : n6374_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6393_o = n6374_o & n6384_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6395_o = n6374_o & n6384_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6396_o = n6374_o & n6384_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6397_o = n6393_o & n6374_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6399_o = n6395_o & n6374_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6400_o = n6396_o & n6374_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6402_o = challenge == 8'b00011100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6403_o = sortie_ro[28];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6404_o = n6415_o ? n6403_o : n6386_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6406_o = n6417_o ? 1'b1 : n6388_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6410_o = n6418_o ? 1'b0 : n6392_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6411_o = n6392_o & n6402_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6413_o = n6392_o & n6402_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6414_o = n6392_o & n6402_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6415_o = n6411_o & n6392_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6417_o = n6413_o & n6392_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6418_o = n6414_o & n6392_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6420_o = challenge == 8'b00011101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6421_o = sortie_ro[29];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6422_o = n6433_o ? n6421_o : n6404_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6424_o = n6435_o ? 1'b1 : n6406_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6428_o = n6436_o ? 1'b0 : n6410_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6429_o = n6410_o & n6420_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6431_o = n6410_o & n6420_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6432_o = n6410_o & n6420_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6433_o = n6429_o & n6410_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6435_o = n6431_o & n6410_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6436_o = n6432_o & n6410_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6438_o = challenge == 8'b00011110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6439_o = sortie_ro[30];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6440_o = n6451_o ? n6439_o : n6422_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6442_o = n6453_o ? 1'b1 : n6424_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6446_o = n6454_o ? 1'b0 : n6428_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6447_o = n6428_o & n6438_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6449_o = n6428_o & n6438_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6450_o = n6428_o & n6438_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6451_o = n6447_o & n6428_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6453_o = n6449_o & n6428_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6454_o = n6450_o & n6428_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6456_o = challenge == 8'b00011111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6457_o = sortie_ro[31];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6458_o = n6469_o ? n6457_o : n6440_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6460_o = n6471_o ? 1'b1 : n6442_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6464_o = n6472_o ? 1'b0 : n6446_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6465_o = n6446_o & n6456_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6467_o = n6446_o & n6456_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6468_o = n6446_o & n6456_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6469_o = n6465_o & n6446_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6471_o = n6467_o & n6446_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6472_o = n6468_o & n6446_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6474_o = challenge == 8'b00100000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6475_o = sortie_ro[32];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6476_o = n6487_o ? n6475_o : n6458_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6478_o = n6489_o ? 1'b1 : n6460_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6482_o = n6490_o ? 1'b0 : n6464_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6483_o = n6464_o & n6474_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6485_o = n6464_o & n6474_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6486_o = n6464_o & n6474_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6487_o = n6483_o & n6464_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6489_o = n6485_o & n6464_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6490_o = n6486_o & n6464_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6492_o = challenge == 8'b00100001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6493_o = sortie_ro[33];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6494_o = n6505_o ? n6493_o : n6476_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6496_o = n6507_o ? 1'b1 : n6478_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6500_o = n6508_o ? 1'b0 : n6482_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6501_o = n6482_o & n6492_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6503_o = n6482_o & n6492_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6504_o = n6482_o & n6492_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6505_o = n6501_o & n6482_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6507_o = n6503_o & n6482_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6508_o = n6504_o & n6482_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6510_o = challenge == 8'b00100010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6511_o = sortie_ro[34];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6512_o = n6523_o ? n6511_o : n6494_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6514_o = n6525_o ? 1'b1 : n6496_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6518_o = n6526_o ? 1'b0 : n6500_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6519_o = n6500_o & n6510_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6521_o = n6500_o & n6510_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6522_o = n6500_o & n6510_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6523_o = n6519_o & n6500_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6525_o = n6521_o & n6500_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6526_o = n6522_o & n6500_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6528_o = challenge == 8'b00100011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6529_o = sortie_ro[35];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6530_o = n6541_o ? n6529_o : n6512_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6532_o = n6543_o ? 1'b1 : n6514_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6536_o = n6544_o ? 1'b0 : n6518_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6537_o = n6518_o & n6528_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6539_o = n6518_o & n6528_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6540_o = n6518_o & n6528_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6541_o = n6537_o & n6518_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6543_o = n6539_o & n6518_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6544_o = n6540_o & n6518_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6546_o = challenge == 8'b00100100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6547_o = sortie_ro[36];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6548_o = n6559_o ? n6547_o : n6530_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6550_o = n6561_o ? 1'b1 : n6532_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6554_o = n6562_o ? 1'b0 : n6536_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6555_o = n6536_o & n6546_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6557_o = n6536_o & n6546_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6558_o = n6536_o & n6546_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6559_o = n6555_o & n6536_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6561_o = n6557_o & n6536_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6562_o = n6558_o & n6536_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6564_o = challenge == 8'b00100101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6565_o = sortie_ro[37];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6566_o = n6577_o ? n6565_o : n6548_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6568_o = n6579_o ? 1'b1 : n6550_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6572_o = n6580_o ? 1'b0 : n6554_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6573_o = n6554_o & n6564_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6575_o = n6554_o & n6564_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6576_o = n6554_o & n6564_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6577_o = n6573_o & n6554_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6579_o = n6575_o & n6554_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6580_o = n6576_o & n6554_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6582_o = challenge == 8'b00100110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6583_o = sortie_ro[38];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6584_o = n6595_o ? n6583_o : n6566_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6586_o = n6597_o ? 1'b1 : n6568_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6590_o = n6598_o ? 1'b0 : n6572_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6591_o = n6572_o & n6582_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6593_o = n6572_o & n6582_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6594_o = n6572_o & n6582_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6595_o = n6591_o & n6572_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6597_o = n6593_o & n6572_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6598_o = n6594_o & n6572_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6600_o = challenge == 8'b00100111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6601_o = sortie_ro[39];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6602_o = n6613_o ? n6601_o : n6584_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6604_o = n6615_o ? 1'b1 : n6586_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6608_o = n6616_o ? 1'b0 : n6590_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6609_o = n6590_o & n6600_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6611_o = n6590_o & n6600_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6612_o = n6590_o & n6600_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6613_o = n6609_o & n6590_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6615_o = n6611_o & n6590_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6616_o = n6612_o & n6590_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6618_o = challenge == 8'b00101000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6619_o = sortie_ro[40];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6620_o = n6631_o ? n6619_o : n6602_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6622_o = n6633_o ? 1'b1 : n6604_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6626_o = n6634_o ? 1'b0 : n6608_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6627_o = n6608_o & n6618_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6629_o = n6608_o & n6618_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6630_o = n6608_o & n6618_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6631_o = n6627_o & n6608_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6633_o = n6629_o & n6608_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6634_o = n6630_o & n6608_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6636_o = challenge == 8'b00101001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6637_o = sortie_ro[41];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6638_o = n6649_o ? n6637_o : n6620_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6640_o = n6651_o ? 1'b1 : n6622_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6644_o = n6652_o ? 1'b0 : n6626_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6645_o = n6626_o & n6636_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6647_o = n6626_o & n6636_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6648_o = n6626_o & n6636_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6649_o = n6645_o & n6626_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6651_o = n6647_o & n6626_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6652_o = n6648_o & n6626_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6654_o = challenge == 8'b00101010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6655_o = sortie_ro[42];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6656_o = n6667_o ? n6655_o : n6638_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6658_o = n6669_o ? 1'b1 : n6640_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6662_o = n6670_o ? 1'b0 : n6644_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6663_o = n6644_o & n6654_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6665_o = n6644_o & n6654_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6666_o = n6644_o & n6654_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6667_o = n6663_o & n6644_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6669_o = n6665_o & n6644_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6670_o = n6666_o & n6644_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6672_o = challenge == 8'b00101011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6673_o = sortie_ro[43];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6674_o = n6685_o ? n6673_o : n6656_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6676_o = n6687_o ? 1'b1 : n6658_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6680_o = n6688_o ? 1'b0 : n6662_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6681_o = n6662_o & n6672_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6683_o = n6662_o & n6672_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6684_o = n6662_o & n6672_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6685_o = n6681_o & n6662_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6687_o = n6683_o & n6662_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6688_o = n6684_o & n6662_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6690_o = challenge == 8'b00101100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6691_o = sortie_ro[44];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6692_o = n6703_o ? n6691_o : n6674_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6694_o = n6705_o ? 1'b1 : n6676_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6698_o = n6706_o ? 1'b0 : n6680_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6699_o = n6680_o & n6690_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6701_o = n6680_o & n6690_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6702_o = n6680_o & n6690_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6703_o = n6699_o & n6680_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6705_o = n6701_o & n6680_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6706_o = n6702_o & n6680_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6708_o = challenge == 8'b00101101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6709_o = sortie_ro[45];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6710_o = n6721_o ? n6709_o : n6692_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6712_o = n6723_o ? 1'b1 : n6694_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6716_o = n6724_o ? 1'b0 : n6698_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6717_o = n6698_o & n6708_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6719_o = n6698_o & n6708_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6720_o = n6698_o & n6708_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6721_o = n6717_o & n6698_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6723_o = n6719_o & n6698_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6724_o = n6720_o & n6698_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6726_o = challenge == 8'b00101110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6727_o = sortie_ro[46];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6728_o = n6739_o ? n6727_o : n6710_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6730_o = n6741_o ? 1'b1 : n6712_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6734_o = n6742_o ? 1'b0 : n6716_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6735_o = n6716_o & n6726_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6737_o = n6716_o & n6726_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6738_o = n6716_o & n6726_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6739_o = n6735_o & n6716_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6741_o = n6737_o & n6716_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6742_o = n6738_o & n6716_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6744_o = challenge == 8'b00101111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6745_o = sortie_ro[47];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6746_o = n6757_o ? n6745_o : n6728_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6748_o = n6759_o ? 1'b1 : n6730_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6752_o = n6760_o ? 1'b0 : n6734_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6753_o = n6734_o & n6744_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6755_o = n6734_o & n6744_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6756_o = n6734_o & n6744_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6757_o = n6753_o & n6734_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6759_o = n6755_o & n6734_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6760_o = n6756_o & n6734_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6762_o = challenge == 8'b00110000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6763_o = sortie_ro[48];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6764_o = n6775_o ? n6763_o : n6746_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6766_o = n6777_o ? 1'b1 : n6748_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6770_o = n6778_o ? 1'b0 : n6752_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6771_o = n6752_o & n6762_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6773_o = n6752_o & n6762_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6774_o = n6752_o & n6762_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6775_o = n6771_o & n6752_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6777_o = n6773_o & n6752_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6778_o = n6774_o & n6752_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6780_o = challenge == 8'b00110001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6781_o = sortie_ro[49];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6782_o = n6793_o ? n6781_o : n6764_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6784_o = n6795_o ? 1'b1 : n6766_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6788_o = n6796_o ? 1'b0 : n6770_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6789_o = n6770_o & n6780_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6791_o = n6770_o & n6780_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6792_o = n6770_o & n6780_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6793_o = n6789_o & n6770_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6795_o = n6791_o & n6770_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6796_o = n6792_o & n6770_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6798_o = challenge == 8'b00110010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6799_o = sortie_ro[50];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6800_o = n6811_o ? n6799_o : n6782_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6802_o = n6813_o ? 1'b1 : n6784_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6806_o = n6814_o ? 1'b0 : n6788_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6807_o = n6788_o & n6798_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6809_o = n6788_o & n6798_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6810_o = n6788_o & n6798_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6811_o = n6807_o & n6788_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6813_o = n6809_o & n6788_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6814_o = n6810_o & n6788_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6816_o = challenge == 8'b00110011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6817_o = sortie_ro[51];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6818_o = n6829_o ? n6817_o : n6800_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6820_o = n6831_o ? 1'b1 : n6802_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6824_o = n6832_o ? 1'b0 : n6806_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6825_o = n6806_o & n6816_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6827_o = n6806_o & n6816_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6828_o = n6806_o & n6816_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6829_o = n6825_o & n6806_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6831_o = n6827_o & n6806_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6832_o = n6828_o & n6806_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6834_o = challenge == 8'b00110100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6835_o = sortie_ro[52];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6836_o = n6847_o ? n6835_o : n6818_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6838_o = n6849_o ? 1'b1 : n6820_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6842_o = n6850_o ? 1'b0 : n6824_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6843_o = n6824_o & n6834_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6845_o = n6824_o & n6834_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6846_o = n6824_o & n6834_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6847_o = n6843_o & n6824_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6849_o = n6845_o & n6824_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6850_o = n6846_o & n6824_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6852_o = challenge == 8'b00110101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6853_o = sortie_ro[53];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6854_o = n6865_o ? n6853_o : n6836_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6856_o = n6867_o ? 1'b1 : n6838_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6860_o = n6868_o ? 1'b0 : n6842_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6861_o = n6842_o & n6852_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6863_o = n6842_o & n6852_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6864_o = n6842_o & n6852_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6865_o = n6861_o & n6842_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6867_o = n6863_o & n6842_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6868_o = n6864_o & n6842_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6870_o = challenge == 8'b00110110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6871_o = sortie_ro[54];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6872_o = n6883_o ? n6871_o : n6854_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6874_o = n6885_o ? 1'b1 : n6856_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6878_o = n6886_o ? 1'b0 : n6860_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6879_o = n6860_o & n6870_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6881_o = n6860_o & n6870_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6882_o = n6860_o & n6870_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6883_o = n6879_o & n6860_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6885_o = n6881_o & n6860_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6886_o = n6882_o & n6860_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6888_o = challenge == 8'b00110111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6889_o = sortie_ro[55];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6890_o = n6901_o ? n6889_o : n6872_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6892_o = n6903_o ? 1'b1 : n6874_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6896_o = n6904_o ? 1'b0 : n6878_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6897_o = n6878_o & n6888_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6899_o = n6878_o & n6888_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6900_o = n6878_o & n6888_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6901_o = n6897_o & n6878_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6903_o = n6899_o & n6878_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6904_o = n6900_o & n6878_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6906_o = challenge == 8'b00111000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6907_o = sortie_ro[56];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6908_o = n6919_o ? n6907_o : n6890_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6910_o = n6921_o ? 1'b1 : n6892_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6914_o = n6922_o ? 1'b0 : n6896_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6915_o = n6896_o & n6906_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6917_o = n6896_o & n6906_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6918_o = n6896_o & n6906_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6919_o = n6915_o & n6896_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6921_o = n6917_o & n6896_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6922_o = n6918_o & n6896_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6924_o = challenge == 8'b00111001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6925_o = sortie_ro[57];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6926_o = n6937_o ? n6925_o : n6908_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6928_o = n6939_o ? 1'b1 : n6910_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6932_o = n6940_o ? 1'b0 : n6914_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6933_o = n6914_o & n6924_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6935_o = n6914_o & n6924_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6936_o = n6914_o & n6924_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6937_o = n6933_o & n6914_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6939_o = n6935_o & n6914_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6940_o = n6936_o & n6914_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6942_o = challenge == 8'b00111010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6943_o = sortie_ro[58];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6944_o = n6955_o ? n6943_o : n6926_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6946_o = n6957_o ? 1'b1 : n6928_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6950_o = n6958_o ? 1'b0 : n6932_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6951_o = n6932_o & n6942_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6953_o = n6932_o & n6942_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6954_o = n6932_o & n6942_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6955_o = n6951_o & n6932_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6957_o = n6953_o & n6932_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6958_o = n6954_o & n6932_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6960_o = challenge == 8'b00111011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6961_o = sortie_ro[59];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6962_o = n6973_o ? n6961_o : n6944_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6964_o = n6975_o ? 1'b1 : n6946_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6968_o = n6976_o ? 1'b0 : n6950_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6969_o = n6950_o & n6960_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6971_o = n6950_o & n6960_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6972_o = n6950_o & n6960_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6973_o = n6969_o & n6950_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6975_o = n6971_o & n6950_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6976_o = n6972_o & n6950_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6978_o = challenge == 8'b00111100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6979_o = sortie_ro[60];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6980_o = n6991_o ? n6979_o : n6962_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6982_o = n6993_o ? 1'b1 : n6964_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6986_o = n6994_o ? 1'b0 : n6968_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6987_o = n6968_o & n6978_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6989_o = n6968_o & n6978_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6990_o = n6968_o & n6978_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6991_o = n6987_o & n6968_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6993_o = n6989_o & n6968_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6994_o = n6990_o & n6968_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n6996_o = challenge == 8'b00111101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n6997_o = sortie_ro[61];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n6998_o = n7009_o ? n6997_o : n6980_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7000_o = n7011_o ? 1'b1 : n6982_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7004_o = n7012_o ? 1'b0 : n6986_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7005_o = n6986_o & n6996_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7007_o = n6986_o & n6996_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7008_o = n6986_o & n6996_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7009_o = n7005_o & n6986_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7011_o = n7007_o & n6986_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7012_o = n7008_o & n6986_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7014_o = challenge == 8'b00111110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7015_o = sortie_ro[62];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7016_o = n7027_o ? n7015_o : n6998_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7018_o = n7029_o ? 1'b1 : n7000_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7022_o = n7030_o ? 1'b0 : n7004_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7023_o = n7004_o & n7014_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7025_o = n7004_o & n7014_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7026_o = n7004_o & n7014_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7027_o = n7023_o & n7004_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7029_o = n7025_o & n7004_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7030_o = n7026_o & n7004_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7032_o = challenge == 8'b00111111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7033_o = sortie_ro[63];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7034_o = n7045_o ? n7033_o : n7016_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7036_o = n7047_o ? 1'b1 : n7018_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7040_o = n7048_o ? 1'b0 : n7022_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7041_o = n7022_o & n7032_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7043_o = n7022_o & n7032_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7044_o = n7022_o & n7032_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7045_o = n7041_o & n7022_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7047_o = n7043_o & n7022_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7048_o = n7044_o & n7022_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7050_o = challenge == 8'b01000000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7051_o = sortie_ro[64];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7052_o = n7063_o ? n7051_o : n7034_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7054_o = n7065_o ? 1'b1 : n7036_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7058_o = n7066_o ? 1'b0 : n7040_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7059_o = n7040_o & n7050_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7061_o = n7040_o & n7050_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7062_o = n7040_o & n7050_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7063_o = n7059_o & n7040_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7065_o = n7061_o & n7040_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7066_o = n7062_o & n7040_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7068_o = challenge == 8'b01000001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7069_o = sortie_ro[65];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7070_o = n7081_o ? n7069_o : n7052_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7072_o = n7083_o ? 1'b1 : n7054_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7076_o = n7084_o ? 1'b0 : n7058_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7077_o = n7058_o & n7068_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7079_o = n7058_o & n7068_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7080_o = n7058_o & n7068_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7081_o = n7077_o & n7058_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7083_o = n7079_o & n7058_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7084_o = n7080_o & n7058_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7086_o = challenge == 8'b01000010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7087_o = sortie_ro[66];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7088_o = n7099_o ? n7087_o : n7070_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7090_o = n7101_o ? 1'b1 : n7072_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7094_o = n7102_o ? 1'b0 : n7076_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7095_o = n7076_o & n7086_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7097_o = n7076_o & n7086_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7098_o = n7076_o & n7086_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7099_o = n7095_o & n7076_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7101_o = n7097_o & n7076_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7102_o = n7098_o & n7076_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7104_o = challenge == 8'b01000011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7105_o = sortie_ro[67];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7106_o = n7117_o ? n7105_o : n7088_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7108_o = n7119_o ? 1'b1 : n7090_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7112_o = n7120_o ? 1'b0 : n7094_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7113_o = n7094_o & n7104_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7115_o = n7094_o & n7104_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7116_o = n7094_o & n7104_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7117_o = n7113_o & n7094_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7119_o = n7115_o & n7094_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7120_o = n7116_o & n7094_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7122_o = challenge == 8'b01000100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7123_o = sortie_ro[68];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7124_o = n7135_o ? n7123_o : n7106_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7126_o = n7137_o ? 1'b1 : n7108_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7130_o = n7138_o ? 1'b0 : n7112_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7131_o = n7112_o & n7122_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7133_o = n7112_o & n7122_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7134_o = n7112_o & n7122_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7135_o = n7131_o & n7112_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7137_o = n7133_o & n7112_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7138_o = n7134_o & n7112_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7140_o = challenge == 8'b01000101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7141_o = sortie_ro[69];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7142_o = n7153_o ? n7141_o : n7124_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7144_o = n7155_o ? 1'b1 : n7126_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7148_o = n7156_o ? 1'b0 : n7130_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7149_o = n7130_o & n7140_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7151_o = n7130_o & n7140_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7152_o = n7130_o & n7140_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7153_o = n7149_o & n7130_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7155_o = n7151_o & n7130_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7156_o = n7152_o & n7130_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7158_o = challenge == 8'b01000110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7159_o = sortie_ro[70];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7160_o = n7171_o ? n7159_o : n7142_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7162_o = n7173_o ? 1'b1 : n7144_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7166_o = n7174_o ? 1'b0 : n7148_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7167_o = n7148_o & n7158_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7169_o = n7148_o & n7158_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7170_o = n7148_o & n7158_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7171_o = n7167_o & n7148_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7173_o = n7169_o & n7148_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7174_o = n7170_o & n7148_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7176_o = challenge == 8'b01000111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7177_o = sortie_ro[71];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7178_o = n7189_o ? n7177_o : n7160_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7180_o = n7191_o ? 1'b1 : n7162_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7184_o = n7192_o ? 1'b0 : n7166_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7185_o = n7166_o & n7176_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7187_o = n7166_o & n7176_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7188_o = n7166_o & n7176_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7189_o = n7185_o & n7166_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7191_o = n7187_o & n7166_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7192_o = n7188_o & n7166_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7194_o = challenge == 8'b01001000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7195_o = sortie_ro[72];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7196_o = n7207_o ? n7195_o : n7178_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7198_o = n7209_o ? 1'b1 : n7180_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7202_o = n7210_o ? 1'b0 : n7184_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7203_o = n7184_o & n7194_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7205_o = n7184_o & n7194_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7206_o = n7184_o & n7194_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7207_o = n7203_o & n7184_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7209_o = n7205_o & n7184_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7210_o = n7206_o & n7184_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7212_o = challenge == 8'b01001001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7213_o = sortie_ro[73];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7214_o = n7225_o ? n7213_o : n7196_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7216_o = n7227_o ? 1'b1 : n7198_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7220_o = n7228_o ? 1'b0 : n7202_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7221_o = n7202_o & n7212_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7223_o = n7202_o & n7212_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7224_o = n7202_o & n7212_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7225_o = n7221_o & n7202_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7227_o = n7223_o & n7202_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7228_o = n7224_o & n7202_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7230_o = challenge == 8'b01001010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7231_o = sortie_ro[74];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7232_o = n7243_o ? n7231_o : n7214_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7234_o = n7245_o ? 1'b1 : n7216_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7238_o = n7246_o ? 1'b0 : n7220_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7239_o = n7220_o & n7230_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7241_o = n7220_o & n7230_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7242_o = n7220_o & n7230_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7243_o = n7239_o & n7220_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7245_o = n7241_o & n7220_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7246_o = n7242_o & n7220_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7248_o = challenge == 8'b01001011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7249_o = sortie_ro[75];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7250_o = n7261_o ? n7249_o : n7232_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7252_o = n7263_o ? 1'b1 : n7234_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7256_o = n7264_o ? 1'b0 : n7238_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7257_o = n7238_o & n7248_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7259_o = n7238_o & n7248_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7260_o = n7238_o & n7248_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7261_o = n7257_o & n7238_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7263_o = n7259_o & n7238_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7264_o = n7260_o & n7238_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7266_o = challenge == 8'b01001100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7267_o = sortie_ro[76];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7268_o = n7279_o ? n7267_o : n7250_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7270_o = n7281_o ? 1'b1 : n7252_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7274_o = n7282_o ? 1'b0 : n7256_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7275_o = n7256_o & n7266_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7277_o = n7256_o & n7266_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7278_o = n7256_o & n7266_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7279_o = n7275_o & n7256_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7281_o = n7277_o & n7256_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7282_o = n7278_o & n7256_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7284_o = challenge == 8'b01001101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7285_o = sortie_ro[77];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7286_o = n7297_o ? n7285_o : n7268_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7288_o = n7299_o ? 1'b1 : n7270_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7292_o = n7300_o ? 1'b0 : n7274_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7293_o = n7274_o & n7284_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7295_o = n7274_o & n7284_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7296_o = n7274_o & n7284_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7297_o = n7293_o & n7274_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7299_o = n7295_o & n7274_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7300_o = n7296_o & n7274_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7302_o = challenge == 8'b01001110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7303_o = sortie_ro[78];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7304_o = n7315_o ? n7303_o : n7286_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7306_o = n7317_o ? 1'b1 : n7288_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7310_o = n7318_o ? 1'b0 : n7292_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7311_o = n7292_o & n7302_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7313_o = n7292_o & n7302_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7314_o = n7292_o & n7302_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7315_o = n7311_o & n7292_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7317_o = n7313_o & n7292_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7318_o = n7314_o & n7292_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7320_o = challenge == 8'b01001111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7321_o = sortie_ro[79];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7322_o = n7333_o ? n7321_o : n7304_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7324_o = n7335_o ? 1'b1 : n7306_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7328_o = n7336_o ? 1'b0 : n7310_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7329_o = n7310_o & n7320_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7331_o = n7310_o & n7320_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7332_o = n7310_o & n7320_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7333_o = n7329_o & n7310_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7335_o = n7331_o & n7310_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7336_o = n7332_o & n7310_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7338_o = challenge == 8'b01010000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7339_o = sortie_ro[80];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7340_o = n7351_o ? n7339_o : n7322_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7342_o = n7353_o ? 1'b1 : n7324_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7346_o = n7354_o ? 1'b0 : n7328_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7347_o = n7328_o & n7338_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7349_o = n7328_o & n7338_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7350_o = n7328_o & n7338_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7351_o = n7347_o & n7328_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7353_o = n7349_o & n7328_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7354_o = n7350_o & n7328_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7356_o = challenge == 8'b01010001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7357_o = sortie_ro[81];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7358_o = n7369_o ? n7357_o : n7340_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7360_o = n7371_o ? 1'b1 : n7342_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7364_o = n7372_o ? 1'b0 : n7346_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7365_o = n7346_o & n7356_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7367_o = n7346_o & n7356_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7368_o = n7346_o & n7356_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7369_o = n7365_o & n7346_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7371_o = n7367_o & n7346_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7372_o = n7368_o & n7346_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7374_o = challenge == 8'b01010010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7375_o = sortie_ro[82];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7376_o = n7387_o ? n7375_o : n7358_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7378_o = n7389_o ? 1'b1 : n7360_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7382_o = n7390_o ? 1'b0 : n7364_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7383_o = n7364_o & n7374_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7385_o = n7364_o & n7374_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7386_o = n7364_o & n7374_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7387_o = n7383_o & n7364_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7389_o = n7385_o & n7364_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7390_o = n7386_o & n7364_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7392_o = challenge == 8'b01010011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7393_o = sortie_ro[83];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7394_o = n7405_o ? n7393_o : n7376_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7396_o = n7407_o ? 1'b1 : n7378_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7400_o = n7408_o ? 1'b0 : n7382_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7401_o = n7382_o & n7392_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7403_o = n7382_o & n7392_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7404_o = n7382_o & n7392_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7405_o = n7401_o & n7382_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7407_o = n7403_o & n7382_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7408_o = n7404_o & n7382_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7410_o = challenge == 8'b01010100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7411_o = sortie_ro[84];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7412_o = n7423_o ? n7411_o : n7394_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7414_o = n7425_o ? 1'b1 : n7396_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7418_o = n7426_o ? 1'b0 : n7400_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7419_o = n7400_o & n7410_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7421_o = n7400_o & n7410_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7422_o = n7400_o & n7410_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7423_o = n7419_o & n7400_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7425_o = n7421_o & n7400_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7426_o = n7422_o & n7400_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7428_o = challenge == 8'b01010101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7429_o = sortie_ro[85];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7430_o = n7441_o ? n7429_o : n7412_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7432_o = n7443_o ? 1'b1 : n7414_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7436_o = n7444_o ? 1'b0 : n7418_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7437_o = n7418_o & n7428_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7439_o = n7418_o & n7428_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7440_o = n7418_o & n7428_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7441_o = n7437_o & n7418_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7443_o = n7439_o & n7418_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7444_o = n7440_o & n7418_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7446_o = challenge == 8'b01010110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7447_o = sortie_ro[86];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7448_o = n7459_o ? n7447_o : n7430_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7450_o = n7461_o ? 1'b1 : n7432_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7454_o = n7462_o ? 1'b0 : n7436_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7455_o = n7436_o & n7446_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7457_o = n7436_o & n7446_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7458_o = n7436_o & n7446_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7459_o = n7455_o & n7436_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7461_o = n7457_o & n7436_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7462_o = n7458_o & n7436_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7464_o = challenge == 8'b01010111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7465_o = sortie_ro[87];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7466_o = n7477_o ? n7465_o : n7448_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7468_o = n7479_o ? 1'b1 : n7450_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7472_o = n7480_o ? 1'b0 : n7454_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7473_o = n7454_o & n7464_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7475_o = n7454_o & n7464_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7476_o = n7454_o & n7464_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7477_o = n7473_o & n7454_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7479_o = n7475_o & n7454_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7480_o = n7476_o & n7454_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7482_o = challenge == 8'b01011000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7483_o = sortie_ro[88];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7484_o = n7495_o ? n7483_o : n7466_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7486_o = n7497_o ? 1'b1 : n7468_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7490_o = n7498_o ? 1'b0 : n7472_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7491_o = n7472_o & n7482_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7493_o = n7472_o & n7482_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7494_o = n7472_o & n7482_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7495_o = n7491_o & n7472_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7497_o = n7493_o & n7472_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7498_o = n7494_o & n7472_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7500_o = challenge == 8'b01011001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7501_o = sortie_ro[89];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7502_o = n7513_o ? n7501_o : n7484_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7504_o = n7515_o ? 1'b1 : n7486_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7508_o = n7516_o ? 1'b0 : n7490_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7509_o = n7490_o & n7500_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7511_o = n7490_o & n7500_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7512_o = n7490_o & n7500_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7513_o = n7509_o & n7490_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7515_o = n7511_o & n7490_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7516_o = n7512_o & n7490_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7518_o = challenge == 8'b01011010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7519_o = sortie_ro[90];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7520_o = n7531_o ? n7519_o : n7502_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7522_o = n7533_o ? 1'b1 : n7504_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7526_o = n7534_o ? 1'b0 : n7508_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7527_o = n7508_o & n7518_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7529_o = n7508_o & n7518_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7530_o = n7508_o & n7518_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7531_o = n7527_o & n7508_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7533_o = n7529_o & n7508_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7534_o = n7530_o & n7508_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7536_o = challenge == 8'b01011011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7537_o = sortie_ro[91];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7538_o = n7549_o ? n7537_o : n7520_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7540_o = n7551_o ? 1'b1 : n7522_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7544_o = n7552_o ? 1'b0 : n7526_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7545_o = n7526_o & n7536_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7547_o = n7526_o & n7536_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7548_o = n7526_o & n7536_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7549_o = n7545_o & n7526_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7551_o = n7547_o & n7526_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7552_o = n7548_o & n7526_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7554_o = challenge == 8'b01011100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7555_o = sortie_ro[92];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7556_o = n7567_o ? n7555_o : n7538_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7558_o = n7569_o ? 1'b1 : n7540_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7562_o = n7570_o ? 1'b0 : n7544_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7563_o = n7544_o & n7554_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7565_o = n7544_o & n7554_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7566_o = n7544_o & n7554_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7567_o = n7563_o & n7544_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7569_o = n7565_o & n7544_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7570_o = n7566_o & n7544_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7572_o = challenge == 8'b01011101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7573_o = sortie_ro[93];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7574_o = n7585_o ? n7573_o : n7556_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7576_o = n7587_o ? 1'b1 : n7558_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7580_o = n7588_o ? 1'b0 : n7562_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7581_o = n7562_o & n7572_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7583_o = n7562_o & n7572_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7584_o = n7562_o & n7572_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7585_o = n7581_o & n7562_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7587_o = n7583_o & n7562_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7588_o = n7584_o & n7562_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7590_o = challenge == 8'b01011110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7591_o = sortie_ro[94];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7592_o = n7603_o ? n7591_o : n7574_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7594_o = n7605_o ? 1'b1 : n7576_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7598_o = n7606_o ? 1'b0 : n7580_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7599_o = n7580_o & n7590_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7601_o = n7580_o & n7590_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7602_o = n7580_o & n7590_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7603_o = n7599_o & n7580_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7605_o = n7601_o & n7580_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7606_o = n7602_o & n7580_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7608_o = challenge == 8'b01011111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7609_o = sortie_ro[95];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7610_o = n7621_o ? n7609_o : n7592_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7612_o = n7623_o ? 1'b1 : n7594_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7616_o = n7624_o ? 1'b0 : n7598_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7617_o = n7598_o & n7608_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7619_o = n7598_o & n7608_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7620_o = n7598_o & n7608_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7621_o = n7617_o & n7598_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7623_o = n7619_o & n7598_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7624_o = n7620_o & n7598_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7626_o = challenge == 8'b01100000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7627_o = sortie_ro[96];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7628_o = n7639_o ? n7627_o : n7610_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7630_o = n7641_o ? 1'b1 : n7612_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7634_o = n7642_o ? 1'b0 : n7616_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7635_o = n7616_o & n7626_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7637_o = n7616_o & n7626_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7638_o = n7616_o & n7626_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7639_o = n7635_o & n7616_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7641_o = n7637_o & n7616_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7642_o = n7638_o & n7616_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7644_o = challenge == 8'b01100001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7645_o = sortie_ro[97];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7646_o = n7657_o ? n7645_o : n7628_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7648_o = n7659_o ? 1'b1 : n7630_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7652_o = n7660_o ? 1'b0 : n7634_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7653_o = n7634_o & n7644_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7655_o = n7634_o & n7644_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7656_o = n7634_o & n7644_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7657_o = n7653_o & n7634_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7659_o = n7655_o & n7634_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7660_o = n7656_o & n7634_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7662_o = challenge == 8'b01100010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7663_o = sortie_ro[98];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7664_o = n7675_o ? n7663_o : n7646_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7666_o = n7677_o ? 1'b1 : n7648_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7670_o = n7678_o ? 1'b0 : n7652_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7671_o = n7652_o & n7662_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7673_o = n7652_o & n7662_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7674_o = n7652_o & n7662_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7675_o = n7671_o & n7652_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7677_o = n7673_o & n7652_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7678_o = n7674_o & n7652_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7680_o = challenge == 8'b01100011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7681_o = sortie_ro[99];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7682_o = n7693_o ? n7681_o : n7664_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7684_o = n7695_o ? 1'b1 : n7666_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7688_o = n7696_o ? 1'b0 : n7670_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7689_o = n7670_o & n7680_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7691_o = n7670_o & n7680_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7692_o = n7670_o & n7680_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7693_o = n7689_o & n7670_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7695_o = n7691_o & n7670_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7696_o = n7692_o & n7670_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7698_o = challenge == 8'b01100100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7699_o = sortie_ro[100];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7700_o = n7711_o ? n7699_o : n7682_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7702_o = n7713_o ? 1'b1 : n7684_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7706_o = n7714_o ? 1'b0 : n7688_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7707_o = n7688_o & n7698_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7709_o = n7688_o & n7698_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7710_o = n7688_o & n7698_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7711_o = n7707_o & n7688_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7713_o = n7709_o & n7688_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7714_o = n7710_o & n7688_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7716_o = challenge == 8'b01100101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7717_o = sortie_ro[101];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7718_o = n7729_o ? n7717_o : n7700_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7720_o = n7731_o ? 1'b1 : n7702_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7724_o = n7732_o ? 1'b0 : n7706_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7725_o = n7706_o & n7716_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7727_o = n7706_o & n7716_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7728_o = n7706_o & n7716_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7729_o = n7725_o & n7706_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7731_o = n7727_o & n7706_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7732_o = n7728_o & n7706_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7734_o = challenge == 8'b01100110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7735_o = sortie_ro[102];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7736_o = n7747_o ? n7735_o : n7718_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7738_o = n7749_o ? 1'b1 : n7720_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7742_o = n7750_o ? 1'b0 : n7724_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7743_o = n7724_o & n7734_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7745_o = n7724_o & n7734_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7746_o = n7724_o & n7734_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7747_o = n7743_o & n7724_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7749_o = n7745_o & n7724_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7750_o = n7746_o & n7724_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7752_o = challenge == 8'b01100111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7753_o = sortie_ro[103];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7754_o = n7765_o ? n7753_o : n7736_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7756_o = n7767_o ? 1'b1 : n7738_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7760_o = n7768_o ? 1'b0 : n7742_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7761_o = n7742_o & n7752_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7763_o = n7742_o & n7752_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7764_o = n7742_o & n7752_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7765_o = n7761_o & n7742_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7767_o = n7763_o & n7742_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7768_o = n7764_o & n7742_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7770_o = challenge == 8'b01101000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7771_o = sortie_ro[104];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7772_o = n7783_o ? n7771_o : n7754_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7774_o = n7785_o ? 1'b1 : n7756_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7778_o = n7786_o ? 1'b0 : n7760_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7779_o = n7760_o & n7770_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7781_o = n7760_o & n7770_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7782_o = n7760_o & n7770_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7783_o = n7779_o & n7760_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7785_o = n7781_o & n7760_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7786_o = n7782_o & n7760_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7788_o = challenge == 8'b01101001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7789_o = sortie_ro[105];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7790_o = n7801_o ? n7789_o : n7772_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7792_o = n7803_o ? 1'b1 : n7774_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7796_o = n7804_o ? 1'b0 : n7778_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7797_o = n7778_o & n7788_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7799_o = n7778_o & n7788_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7800_o = n7778_o & n7788_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7801_o = n7797_o & n7778_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7803_o = n7799_o & n7778_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7804_o = n7800_o & n7778_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7806_o = challenge == 8'b01101010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7807_o = sortie_ro[106];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7808_o = n7819_o ? n7807_o : n7790_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7810_o = n7821_o ? 1'b1 : n7792_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7814_o = n7822_o ? 1'b0 : n7796_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7815_o = n7796_o & n7806_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7817_o = n7796_o & n7806_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7818_o = n7796_o & n7806_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7819_o = n7815_o & n7796_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7821_o = n7817_o & n7796_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7822_o = n7818_o & n7796_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7824_o = challenge == 8'b01101011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7825_o = sortie_ro[107];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7826_o = n7837_o ? n7825_o : n7808_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7828_o = n7839_o ? 1'b1 : n7810_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7832_o = n7840_o ? 1'b0 : n7814_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7833_o = n7814_o & n7824_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7835_o = n7814_o & n7824_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7836_o = n7814_o & n7824_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7837_o = n7833_o & n7814_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7839_o = n7835_o & n7814_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7840_o = n7836_o & n7814_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7842_o = challenge == 8'b01101100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7843_o = sortie_ro[108];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7844_o = n7855_o ? n7843_o : n7826_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7846_o = n7857_o ? 1'b1 : n7828_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7850_o = n7858_o ? 1'b0 : n7832_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7851_o = n7832_o & n7842_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7853_o = n7832_o & n7842_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7854_o = n7832_o & n7842_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7855_o = n7851_o & n7832_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7857_o = n7853_o & n7832_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7858_o = n7854_o & n7832_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7860_o = challenge == 8'b01101101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7861_o = sortie_ro[109];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7862_o = n7873_o ? n7861_o : n7844_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7864_o = n7875_o ? 1'b1 : n7846_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7868_o = n7876_o ? 1'b0 : n7850_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7869_o = n7850_o & n7860_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7871_o = n7850_o & n7860_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7872_o = n7850_o & n7860_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7873_o = n7869_o & n7850_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7875_o = n7871_o & n7850_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7876_o = n7872_o & n7850_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7878_o = challenge == 8'b01101110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7879_o = sortie_ro[110];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7880_o = n7891_o ? n7879_o : n7862_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7882_o = n7893_o ? 1'b1 : n7864_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7886_o = n7894_o ? 1'b0 : n7868_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7887_o = n7868_o & n7878_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7889_o = n7868_o & n7878_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7890_o = n7868_o & n7878_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7891_o = n7887_o & n7868_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7893_o = n7889_o & n7868_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7894_o = n7890_o & n7868_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7896_o = challenge == 8'b01101111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7897_o = sortie_ro[111];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7898_o = n7909_o ? n7897_o : n7880_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7900_o = n7911_o ? 1'b1 : n7882_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7904_o = n7912_o ? 1'b0 : n7886_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7905_o = n7886_o & n7896_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7907_o = n7886_o & n7896_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7908_o = n7886_o & n7896_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7909_o = n7905_o & n7886_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7911_o = n7907_o & n7886_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7912_o = n7908_o & n7886_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7914_o = challenge == 8'b01110000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7915_o = sortie_ro[112];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7916_o = n7927_o ? n7915_o : n7898_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7918_o = n7929_o ? 1'b1 : n7900_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7922_o = n7930_o ? 1'b0 : n7904_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7923_o = n7904_o & n7914_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7925_o = n7904_o & n7914_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7926_o = n7904_o & n7914_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7927_o = n7923_o & n7904_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7929_o = n7925_o & n7904_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7930_o = n7926_o & n7904_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7932_o = challenge == 8'b01110001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7933_o = sortie_ro[113];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7934_o = n7945_o ? n7933_o : n7916_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7936_o = n7947_o ? 1'b1 : n7918_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7940_o = n7948_o ? 1'b0 : n7922_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7941_o = n7922_o & n7932_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7943_o = n7922_o & n7932_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7944_o = n7922_o & n7932_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7945_o = n7941_o & n7922_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7947_o = n7943_o & n7922_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7948_o = n7944_o & n7922_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7950_o = challenge == 8'b01110010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7951_o = sortie_ro[114];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7952_o = n7963_o ? n7951_o : n7934_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7954_o = n7965_o ? 1'b1 : n7936_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7958_o = n7966_o ? 1'b0 : n7940_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7959_o = n7940_o & n7950_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7961_o = n7940_o & n7950_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7962_o = n7940_o & n7950_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7963_o = n7959_o & n7940_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7965_o = n7961_o & n7940_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7966_o = n7962_o & n7940_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7968_o = challenge == 8'b01110011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7969_o = sortie_ro[115];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7970_o = n7981_o ? n7969_o : n7952_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7972_o = n7983_o ? 1'b1 : n7954_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7976_o = n7984_o ? 1'b0 : n7958_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7977_o = n7958_o & n7968_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7979_o = n7958_o & n7968_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7980_o = n7958_o & n7968_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7981_o = n7977_o & n7958_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7983_o = n7979_o & n7958_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7984_o = n7980_o & n7958_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n7986_o = challenge == 8'b01110100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n7987_o = sortie_ro[116];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7988_o = n7999_o ? n7987_o : n7970_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7990_o = n8001_o ? 1'b1 : n7972_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7994_o = n8002_o ? 1'b0 : n7976_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7995_o = n7976_o & n7986_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7997_o = n7976_o & n7986_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7998_o = n7976_o & n7986_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n7999_o = n7995_o & n7976_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8001_o = n7997_o & n7976_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8002_o = n7998_o & n7976_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8004_o = challenge == 8'b01110101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8005_o = sortie_ro[117];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8006_o = n8017_o ? n8005_o : n7988_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8008_o = n8019_o ? 1'b1 : n7990_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8012_o = n8020_o ? 1'b0 : n7994_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8013_o = n7994_o & n8004_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8015_o = n7994_o & n8004_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8016_o = n7994_o & n8004_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8017_o = n8013_o & n7994_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8019_o = n8015_o & n7994_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8020_o = n8016_o & n7994_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8022_o = challenge == 8'b01110110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8023_o = sortie_ro[118];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8024_o = n8035_o ? n8023_o : n8006_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8026_o = n8037_o ? 1'b1 : n8008_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8030_o = n8038_o ? 1'b0 : n8012_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8031_o = n8012_o & n8022_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8033_o = n8012_o & n8022_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8034_o = n8012_o & n8022_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8035_o = n8031_o & n8012_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8037_o = n8033_o & n8012_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8038_o = n8034_o & n8012_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8040_o = challenge == 8'b01110111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8041_o = sortie_ro[119];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8042_o = n8053_o ? n8041_o : n8024_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8044_o = n8055_o ? 1'b1 : n8026_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8048_o = n8056_o ? 1'b0 : n8030_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8049_o = n8030_o & n8040_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8051_o = n8030_o & n8040_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8052_o = n8030_o & n8040_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8053_o = n8049_o & n8030_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8055_o = n8051_o & n8030_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8056_o = n8052_o & n8030_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8058_o = challenge == 8'b01111000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8059_o = sortie_ro[120];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8060_o = n8071_o ? n8059_o : n8042_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8062_o = n8073_o ? 1'b1 : n8044_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8066_o = n8074_o ? 1'b0 : n8048_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8067_o = n8048_o & n8058_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8069_o = n8048_o & n8058_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8070_o = n8048_o & n8058_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8071_o = n8067_o & n8048_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8073_o = n8069_o & n8048_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8074_o = n8070_o & n8048_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8076_o = challenge == 8'b01111001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8077_o = sortie_ro[121];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8078_o = n8089_o ? n8077_o : n8060_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8080_o = n8091_o ? 1'b1 : n8062_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8084_o = n8092_o ? 1'b0 : n8066_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8085_o = n8066_o & n8076_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8087_o = n8066_o & n8076_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8088_o = n8066_o & n8076_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8089_o = n8085_o & n8066_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8091_o = n8087_o & n8066_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8092_o = n8088_o & n8066_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8094_o = challenge == 8'b01111010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8095_o = sortie_ro[122];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8096_o = n8107_o ? n8095_o : n8078_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8098_o = n8109_o ? 1'b1 : n8080_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8102_o = n8110_o ? 1'b0 : n8084_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8103_o = n8084_o & n8094_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8105_o = n8084_o & n8094_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8106_o = n8084_o & n8094_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8107_o = n8103_o & n8084_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8109_o = n8105_o & n8084_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8110_o = n8106_o & n8084_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8112_o = challenge == 8'b01111011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8113_o = sortie_ro[123];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8114_o = n8125_o ? n8113_o : n8096_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8116_o = n8127_o ? 1'b1 : n8098_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8120_o = n8128_o ? 1'b0 : n8102_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8121_o = n8102_o & n8112_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8123_o = n8102_o & n8112_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8124_o = n8102_o & n8112_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8125_o = n8121_o & n8102_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8127_o = n8123_o & n8102_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8128_o = n8124_o & n8102_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8130_o = challenge == 8'b01111100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8131_o = sortie_ro[124];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8132_o = n8143_o ? n8131_o : n8114_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8134_o = n8145_o ? 1'b1 : n8116_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8138_o = n8146_o ? 1'b0 : n8120_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8139_o = n8120_o & n8130_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8141_o = n8120_o & n8130_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8142_o = n8120_o & n8130_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8143_o = n8139_o & n8120_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8145_o = n8141_o & n8120_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8146_o = n8142_o & n8120_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8148_o = challenge == 8'b01111101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8149_o = sortie_ro[125];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8150_o = n8161_o ? n8149_o : n8132_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8152_o = n8163_o ? 1'b1 : n8134_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8156_o = n8164_o ? 1'b0 : n8138_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8157_o = n8138_o & n8148_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8159_o = n8138_o & n8148_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8160_o = n8138_o & n8148_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8161_o = n8157_o & n8138_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8163_o = n8159_o & n8138_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8164_o = n8160_o & n8138_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8166_o = challenge == 8'b01111110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8167_o = sortie_ro[126];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8168_o = n8179_o ? n8167_o : n8150_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8170_o = n8181_o ? 1'b1 : n8152_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8174_o = n8182_o ? 1'b0 : n8156_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8175_o = n8156_o & n8166_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8177_o = n8156_o & n8166_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8178_o = n8156_o & n8166_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8179_o = n8175_o & n8156_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8181_o = n8177_o & n8156_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8182_o = n8178_o & n8156_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8184_o = challenge == 8'b01111111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8185_o = sortie_ro[127];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8186_o = n8197_o ? n8185_o : n8168_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8188_o = n8199_o ? 1'b1 : n8170_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8192_o = n8200_o ? 1'b0 : n8174_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8193_o = n8174_o & n8184_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8195_o = n8174_o & n8184_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8196_o = n8174_o & n8184_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8197_o = n8193_o & n8174_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8199_o = n8195_o & n8174_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8200_o = n8196_o & n8174_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8202_o = challenge == 8'b10000000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8203_o = sortie_ro[128];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8204_o = n8215_o ? n8203_o : n8186_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8206_o = n8217_o ? 1'b1 : n8188_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8210_o = n8218_o ? 1'b0 : n8192_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8211_o = n8192_o & n8202_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8213_o = n8192_o & n8202_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8214_o = n8192_o & n8202_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8215_o = n8211_o & n8192_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8217_o = n8213_o & n8192_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8218_o = n8214_o & n8192_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8220_o = challenge == 8'b10000001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8221_o = sortie_ro[129];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8222_o = n8233_o ? n8221_o : n8204_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8224_o = n8235_o ? 1'b1 : n8206_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8228_o = n8236_o ? 1'b0 : n8210_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8229_o = n8210_o & n8220_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8231_o = n8210_o & n8220_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8232_o = n8210_o & n8220_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8233_o = n8229_o & n8210_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8235_o = n8231_o & n8210_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8236_o = n8232_o & n8210_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8238_o = challenge == 8'b10000010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8239_o = sortie_ro[130];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8240_o = n8251_o ? n8239_o : n8222_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8242_o = n8253_o ? 1'b1 : n8224_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8246_o = n8254_o ? 1'b0 : n8228_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8247_o = n8228_o & n8238_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8249_o = n8228_o & n8238_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8250_o = n8228_o & n8238_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8251_o = n8247_o & n8228_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8253_o = n8249_o & n8228_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8254_o = n8250_o & n8228_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8256_o = challenge == 8'b10000011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8257_o = sortie_ro[131];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8258_o = n8269_o ? n8257_o : n8240_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8260_o = n8271_o ? 1'b1 : n8242_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8264_o = n8272_o ? 1'b0 : n8246_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8265_o = n8246_o & n8256_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8267_o = n8246_o & n8256_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8268_o = n8246_o & n8256_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8269_o = n8265_o & n8246_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8271_o = n8267_o & n8246_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8272_o = n8268_o & n8246_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8274_o = challenge == 8'b10000100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8275_o = sortie_ro[132];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8276_o = n8287_o ? n8275_o : n8258_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8278_o = n8289_o ? 1'b1 : n8260_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8282_o = n8290_o ? 1'b0 : n8264_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8283_o = n8264_o & n8274_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8285_o = n8264_o & n8274_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8286_o = n8264_o & n8274_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8287_o = n8283_o & n8264_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8289_o = n8285_o & n8264_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8290_o = n8286_o & n8264_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8292_o = challenge == 8'b10000101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8293_o = sortie_ro[133];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8294_o = n8305_o ? n8293_o : n8276_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8296_o = n8307_o ? 1'b1 : n8278_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8300_o = n8308_o ? 1'b0 : n8282_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8301_o = n8282_o & n8292_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8303_o = n8282_o & n8292_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8304_o = n8282_o & n8292_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8305_o = n8301_o & n8282_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8307_o = n8303_o & n8282_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8308_o = n8304_o & n8282_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8310_o = challenge == 8'b10000110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8311_o = sortie_ro[134];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8312_o = n8323_o ? n8311_o : n8294_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8314_o = n8325_o ? 1'b1 : n8296_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8318_o = n8326_o ? 1'b0 : n8300_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8319_o = n8300_o & n8310_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8321_o = n8300_o & n8310_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8322_o = n8300_o & n8310_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8323_o = n8319_o & n8300_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8325_o = n8321_o & n8300_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8326_o = n8322_o & n8300_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8328_o = challenge == 8'b10000111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8329_o = sortie_ro[135];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8330_o = n8341_o ? n8329_o : n8312_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8332_o = n8343_o ? 1'b1 : n8314_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8336_o = n8344_o ? 1'b0 : n8318_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8337_o = n8318_o & n8328_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8339_o = n8318_o & n8328_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8340_o = n8318_o & n8328_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8341_o = n8337_o & n8318_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8343_o = n8339_o & n8318_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8344_o = n8340_o & n8318_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8346_o = challenge == 8'b10001000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8347_o = sortie_ro[136];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8348_o = n8359_o ? n8347_o : n8330_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8350_o = n8361_o ? 1'b1 : n8332_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8354_o = n8362_o ? 1'b0 : n8336_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8355_o = n8336_o & n8346_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8357_o = n8336_o & n8346_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8358_o = n8336_o & n8346_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8359_o = n8355_o & n8336_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8361_o = n8357_o & n8336_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8362_o = n8358_o & n8336_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8364_o = challenge == 8'b10001001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8365_o = sortie_ro[137];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8366_o = n8377_o ? n8365_o : n8348_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8368_o = n8379_o ? 1'b1 : n8350_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8372_o = n8380_o ? 1'b0 : n8354_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8373_o = n8354_o & n8364_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8375_o = n8354_o & n8364_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8376_o = n8354_o & n8364_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8377_o = n8373_o & n8354_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8379_o = n8375_o & n8354_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8380_o = n8376_o & n8354_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8382_o = challenge == 8'b10001010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8383_o = sortie_ro[138];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8384_o = n8395_o ? n8383_o : n8366_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8386_o = n8397_o ? 1'b1 : n8368_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8390_o = n8398_o ? 1'b0 : n8372_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8391_o = n8372_o & n8382_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8393_o = n8372_o & n8382_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8394_o = n8372_o & n8382_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8395_o = n8391_o & n8372_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8397_o = n8393_o & n8372_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8398_o = n8394_o & n8372_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8400_o = challenge == 8'b10001011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8401_o = sortie_ro[139];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8402_o = n8413_o ? n8401_o : n8384_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8404_o = n8415_o ? 1'b1 : n8386_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8408_o = n8416_o ? 1'b0 : n8390_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8409_o = n8390_o & n8400_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8411_o = n8390_o & n8400_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8412_o = n8390_o & n8400_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8413_o = n8409_o & n8390_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8415_o = n8411_o & n8390_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8416_o = n8412_o & n8390_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8418_o = challenge == 8'b10001100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8419_o = sortie_ro[140];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8420_o = n8431_o ? n8419_o : n8402_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8422_o = n8433_o ? 1'b1 : n8404_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8426_o = n8434_o ? 1'b0 : n8408_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8427_o = n8408_o & n8418_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8429_o = n8408_o & n8418_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8430_o = n8408_o & n8418_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8431_o = n8427_o & n8408_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8433_o = n8429_o & n8408_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8434_o = n8430_o & n8408_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8436_o = challenge == 8'b10001101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8437_o = sortie_ro[141];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8438_o = n8449_o ? n8437_o : n8420_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8440_o = n8451_o ? 1'b1 : n8422_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8444_o = n8452_o ? 1'b0 : n8426_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8445_o = n8426_o & n8436_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8447_o = n8426_o & n8436_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8448_o = n8426_o & n8436_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8449_o = n8445_o & n8426_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8451_o = n8447_o & n8426_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8452_o = n8448_o & n8426_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8454_o = challenge == 8'b10001110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8455_o = sortie_ro[142];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8456_o = n8467_o ? n8455_o : n8438_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8458_o = n8469_o ? 1'b1 : n8440_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8462_o = n8470_o ? 1'b0 : n8444_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8463_o = n8444_o & n8454_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8465_o = n8444_o & n8454_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8466_o = n8444_o & n8454_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8467_o = n8463_o & n8444_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8469_o = n8465_o & n8444_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8470_o = n8466_o & n8444_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8472_o = challenge == 8'b10001111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8473_o = sortie_ro[143];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8474_o = n8485_o ? n8473_o : n8456_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8476_o = n8487_o ? 1'b1 : n8458_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8480_o = n8488_o ? 1'b0 : n8462_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8481_o = n8462_o & n8472_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8483_o = n8462_o & n8472_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8484_o = n8462_o & n8472_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8485_o = n8481_o & n8462_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8487_o = n8483_o & n8462_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8488_o = n8484_o & n8462_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8490_o = challenge == 8'b10010000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8491_o = sortie_ro[144];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8492_o = n8503_o ? n8491_o : n8474_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8494_o = n8505_o ? 1'b1 : n8476_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8498_o = n8506_o ? 1'b0 : n8480_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8499_o = n8480_o & n8490_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8501_o = n8480_o & n8490_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8502_o = n8480_o & n8490_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8503_o = n8499_o & n8480_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8505_o = n8501_o & n8480_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8506_o = n8502_o & n8480_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8508_o = challenge == 8'b10010001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8509_o = sortie_ro[145];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8510_o = n8521_o ? n8509_o : n8492_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8512_o = n8523_o ? 1'b1 : n8494_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8516_o = n8524_o ? 1'b0 : n8498_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8517_o = n8498_o & n8508_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8519_o = n8498_o & n8508_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8520_o = n8498_o & n8508_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8521_o = n8517_o & n8498_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8523_o = n8519_o & n8498_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8524_o = n8520_o & n8498_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8526_o = challenge == 8'b10010010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8527_o = sortie_ro[146];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8528_o = n8539_o ? n8527_o : n8510_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8530_o = n8541_o ? 1'b1 : n8512_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8534_o = n8542_o ? 1'b0 : n8516_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8535_o = n8516_o & n8526_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8537_o = n8516_o & n8526_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8538_o = n8516_o & n8526_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8539_o = n8535_o & n8516_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8541_o = n8537_o & n8516_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8542_o = n8538_o & n8516_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8544_o = challenge == 8'b10010011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8545_o = sortie_ro[147];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8546_o = n8557_o ? n8545_o : n8528_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8548_o = n8559_o ? 1'b1 : n8530_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8552_o = n8560_o ? 1'b0 : n8534_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8553_o = n8534_o & n8544_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8555_o = n8534_o & n8544_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8556_o = n8534_o & n8544_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8557_o = n8553_o & n8534_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8559_o = n8555_o & n8534_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8560_o = n8556_o & n8534_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8562_o = challenge == 8'b10010100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8563_o = sortie_ro[148];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8564_o = n8575_o ? n8563_o : n8546_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8566_o = n8577_o ? 1'b1 : n8548_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8570_o = n8578_o ? 1'b0 : n8552_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8571_o = n8552_o & n8562_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8573_o = n8552_o & n8562_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8574_o = n8552_o & n8562_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8575_o = n8571_o & n8552_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8577_o = n8573_o & n8552_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8578_o = n8574_o & n8552_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8580_o = challenge == 8'b10010101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8581_o = sortie_ro[149];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8582_o = n8593_o ? n8581_o : n8564_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8584_o = n8595_o ? 1'b1 : n8566_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8588_o = n8596_o ? 1'b0 : n8570_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8589_o = n8570_o & n8580_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8591_o = n8570_o & n8580_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8592_o = n8570_o & n8580_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8593_o = n8589_o & n8570_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8595_o = n8591_o & n8570_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8596_o = n8592_o & n8570_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8598_o = challenge == 8'b10010110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8599_o = sortie_ro[150];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8600_o = n8611_o ? n8599_o : n8582_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8602_o = n8613_o ? 1'b1 : n8584_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8606_o = n8614_o ? 1'b0 : n8588_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8607_o = n8588_o & n8598_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8609_o = n8588_o & n8598_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8610_o = n8588_o & n8598_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8611_o = n8607_o & n8588_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8613_o = n8609_o & n8588_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8614_o = n8610_o & n8588_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8616_o = challenge == 8'b10010111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8617_o = sortie_ro[151];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8618_o = n8629_o ? n8617_o : n8600_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8620_o = n8631_o ? 1'b1 : n8602_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8624_o = n8632_o ? 1'b0 : n8606_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8625_o = n8606_o & n8616_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8627_o = n8606_o & n8616_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8628_o = n8606_o & n8616_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8629_o = n8625_o & n8606_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8631_o = n8627_o & n8606_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8632_o = n8628_o & n8606_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8634_o = challenge == 8'b10011000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8635_o = sortie_ro[152];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8636_o = n8647_o ? n8635_o : n8618_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8638_o = n8649_o ? 1'b1 : n8620_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8642_o = n8650_o ? 1'b0 : n8624_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8643_o = n8624_o & n8634_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8645_o = n8624_o & n8634_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8646_o = n8624_o & n8634_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8647_o = n8643_o & n8624_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8649_o = n8645_o & n8624_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8650_o = n8646_o & n8624_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8652_o = challenge == 8'b10011001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8653_o = sortie_ro[153];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8654_o = n8665_o ? n8653_o : n8636_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8656_o = n8667_o ? 1'b1 : n8638_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8660_o = n8668_o ? 1'b0 : n8642_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8661_o = n8642_o & n8652_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8663_o = n8642_o & n8652_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8664_o = n8642_o & n8652_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8665_o = n8661_o & n8642_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8667_o = n8663_o & n8642_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8668_o = n8664_o & n8642_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8670_o = challenge == 8'b10011010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8671_o = sortie_ro[154];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8672_o = n8683_o ? n8671_o : n8654_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8674_o = n8685_o ? 1'b1 : n8656_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8678_o = n8686_o ? 1'b0 : n8660_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8679_o = n8660_o & n8670_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8681_o = n8660_o & n8670_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8682_o = n8660_o & n8670_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8683_o = n8679_o & n8660_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8685_o = n8681_o & n8660_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8686_o = n8682_o & n8660_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8688_o = challenge == 8'b10011011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8689_o = sortie_ro[155];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8690_o = n8701_o ? n8689_o : n8672_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8692_o = n8703_o ? 1'b1 : n8674_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8696_o = n8704_o ? 1'b0 : n8678_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8697_o = n8678_o & n8688_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8699_o = n8678_o & n8688_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8700_o = n8678_o & n8688_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8701_o = n8697_o & n8678_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8703_o = n8699_o & n8678_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8704_o = n8700_o & n8678_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8706_o = challenge == 8'b10011100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8707_o = sortie_ro[156];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8708_o = n8719_o ? n8707_o : n8690_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8710_o = n8721_o ? 1'b1 : n8692_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8714_o = n8722_o ? 1'b0 : n8696_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8715_o = n8696_o & n8706_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8717_o = n8696_o & n8706_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8718_o = n8696_o & n8706_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8719_o = n8715_o & n8696_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8721_o = n8717_o & n8696_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8722_o = n8718_o & n8696_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8724_o = challenge == 8'b10011101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8725_o = sortie_ro[157];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8726_o = n8737_o ? n8725_o : n8708_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8728_o = n8739_o ? 1'b1 : n8710_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8732_o = n8740_o ? 1'b0 : n8714_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8733_o = n8714_o & n8724_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8735_o = n8714_o & n8724_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8736_o = n8714_o & n8724_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8737_o = n8733_o & n8714_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8739_o = n8735_o & n8714_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8740_o = n8736_o & n8714_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8742_o = challenge == 8'b10011110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8743_o = sortie_ro[158];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8744_o = n8755_o ? n8743_o : n8726_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8746_o = n8757_o ? 1'b1 : n8728_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8750_o = n8758_o ? 1'b0 : n8732_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8751_o = n8732_o & n8742_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8753_o = n8732_o & n8742_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8754_o = n8732_o & n8742_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8755_o = n8751_o & n8732_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8757_o = n8753_o & n8732_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8758_o = n8754_o & n8732_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8760_o = challenge == 8'b10011111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8761_o = sortie_ro[159];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8762_o = n8773_o ? n8761_o : n8744_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8764_o = n8775_o ? 1'b1 : n8746_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8768_o = n8776_o ? 1'b0 : n8750_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8769_o = n8750_o & n8760_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8771_o = n8750_o & n8760_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8772_o = n8750_o & n8760_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8773_o = n8769_o & n8750_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8775_o = n8771_o & n8750_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8776_o = n8772_o & n8750_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8778_o = challenge == 8'b10100000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8779_o = sortie_ro[160];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8780_o = n8791_o ? n8779_o : n8762_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8782_o = n8793_o ? 1'b1 : n8764_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8786_o = n8794_o ? 1'b0 : n8768_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8787_o = n8768_o & n8778_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8789_o = n8768_o & n8778_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8790_o = n8768_o & n8778_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8791_o = n8787_o & n8768_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8793_o = n8789_o & n8768_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8794_o = n8790_o & n8768_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8796_o = challenge == 8'b10100001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8797_o = sortie_ro[161];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8798_o = n8809_o ? n8797_o : n8780_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8800_o = n8811_o ? 1'b1 : n8782_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8804_o = n8812_o ? 1'b0 : n8786_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8805_o = n8786_o & n8796_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8807_o = n8786_o & n8796_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8808_o = n8786_o & n8796_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8809_o = n8805_o & n8786_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8811_o = n8807_o & n8786_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8812_o = n8808_o & n8786_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8814_o = challenge == 8'b10100010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8815_o = sortie_ro[162];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8816_o = n8827_o ? n8815_o : n8798_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8818_o = n8829_o ? 1'b1 : n8800_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8822_o = n8830_o ? 1'b0 : n8804_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8823_o = n8804_o & n8814_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8825_o = n8804_o & n8814_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8826_o = n8804_o & n8814_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8827_o = n8823_o & n8804_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8829_o = n8825_o & n8804_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8830_o = n8826_o & n8804_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8832_o = challenge == 8'b10100011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8833_o = sortie_ro[163];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8834_o = n8845_o ? n8833_o : n8816_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8836_o = n8847_o ? 1'b1 : n8818_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8840_o = n8848_o ? 1'b0 : n8822_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8841_o = n8822_o & n8832_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8843_o = n8822_o & n8832_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8844_o = n8822_o & n8832_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8845_o = n8841_o & n8822_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8847_o = n8843_o & n8822_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8848_o = n8844_o & n8822_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8850_o = challenge == 8'b10100100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8851_o = sortie_ro[164];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8852_o = n8863_o ? n8851_o : n8834_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8854_o = n8865_o ? 1'b1 : n8836_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8858_o = n8866_o ? 1'b0 : n8840_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8859_o = n8840_o & n8850_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8861_o = n8840_o & n8850_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8862_o = n8840_o & n8850_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8863_o = n8859_o & n8840_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8865_o = n8861_o & n8840_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8866_o = n8862_o & n8840_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8868_o = challenge == 8'b10100101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8869_o = sortie_ro[165];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8870_o = n8881_o ? n8869_o : n8852_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8872_o = n8883_o ? 1'b1 : n8854_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8876_o = n8884_o ? 1'b0 : n8858_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8877_o = n8858_o & n8868_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8879_o = n8858_o & n8868_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8880_o = n8858_o & n8868_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8881_o = n8877_o & n8858_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8883_o = n8879_o & n8858_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8884_o = n8880_o & n8858_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8886_o = challenge == 8'b10100110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8887_o = sortie_ro[166];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8888_o = n8899_o ? n8887_o : n8870_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8890_o = n8901_o ? 1'b1 : n8872_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8894_o = n8902_o ? 1'b0 : n8876_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8895_o = n8876_o & n8886_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8897_o = n8876_o & n8886_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8898_o = n8876_o & n8886_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8899_o = n8895_o & n8876_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8901_o = n8897_o & n8876_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8902_o = n8898_o & n8876_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8904_o = challenge == 8'b10100111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8905_o = sortie_ro[167];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8906_o = n8917_o ? n8905_o : n8888_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8908_o = n8919_o ? 1'b1 : n8890_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8912_o = n8920_o ? 1'b0 : n8894_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8913_o = n8894_o & n8904_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8915_o = n8894_o & n8904_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8916_o = n8894_o & n8904_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8917_o = n8913_o & n8894_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8919_o = n8915_o & n8894_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8920_o = n8916_o & n8894_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8922_o = challenge == 8'b10101000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8923_o = sortie_ro[168];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8924_o = n8935_o ? n8923_o : n8906_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8926_o = n8937_o ? 1'b1 : n8908_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8930_o = n8938_o ? 1'b0 : n8912_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8931_o = n8912_o & n8922_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8933_o = n8912_o & n8922_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8934_o = n8912_o & n8922_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8935_o = n8931_o & n8912_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8937_o = n8933_o & n8912_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8938_o = n8934_o & n8912_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8940_o = challenge == 8'b10101001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8941_o = sortie_ro[169];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8942_o = n8953_o ? n8941_o : n8924_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8944_o = n8955_o ? 1'b1 : n8926_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8948_o = n8956_o ? 1'b0 : n8930_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8949_o = n8930_o & n8940_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8951_o = n8930_o & n8940_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8952_o = n8930_o & n8940_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8953_o = n8949_o & n8930_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8955_o = n8951_o & n8930_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8956_o = n8952_o & n8930_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8958_o = challenge == 8'b10101010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8959_o = sortie_ro[170];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8960_o = n8971_o ? n8959_o : n8942_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8962_o = n8973_o ? 1'b1 : n8944_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8966_o = n8974_o ? 1'b0 : n8948_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8967_o = n8948_o & n8958_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8969_o = n8948_o & n8958_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8970_o = n8948_o & n8958_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8971_o = n8967_o & n8948_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8973_o = n8969_o & n8948_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8974_o = n8970_o & n8948_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8976_o = challenge == 8'b10101011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8977_o = sortie_ro[171];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8978_o = n8989_o ? n8977_o : n8960_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8980_o = n8991_o ? 1'b1 : n8962_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8984_o = n8992_o ? 1'b0 : n8966_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8985_o = n8966_o & n8976_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8987_o = n8966_o & n8976_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8988_o = n8966_o & n8976_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8989_o = n8985_o & n8966_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8991_o = n8987_o & n8966_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8992_o = n8988_o & n8966_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n8994_o = challenge == 8'b10101100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n8995_o = sortie_ro[172];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8996_o = n9007_o ? n8995_o : n8978_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n8998_o = n9009_o ? 1'b1 : n8980_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9002_o = n9010_o ? 1'b0 : n8984_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9003_o = n8984_o & n8994_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9005_o = n8984_o & n8994_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9006_o = n8984_o & n8994_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9007_o = n9003_o & n8984_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9009_o = n9005_o & n8984_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9010_o = n9006_o & n8984_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9012_o = challenge == 8'b10101101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9013_o = sortie_ro[173];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9014_o = n9025_o ? n9013_o : n8996_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9016_o = n9027_o ? 1'b1 : n8998_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9020_o = n9028_o ? 1'b0 : n9002_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9021_o = n9002_o & n9012_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9023_o = n9002_o & n9012_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9024_o = n9002_o & n9012_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9025_o = n9021_o & n9002_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9027_o = n9023_o & n9002_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9028_o = n9024_o & n9002_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9030_o = challenge == 8'b10101110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9031_o = sortie_ro[174];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9032_o = n9043_o ? n9031_o : n9014_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9034_o = n9045_o ? 1'b1 : n9016_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9038_o = n9046_o ? 1'b0 : n9020_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9039_o = n9020_o & n9030_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9041_o = n9020_o & n9030_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9042_o = n9020_o & n9030_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9043_o = n9039_o & n9020_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9045_o = n9041_o & n9020_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9046_o = n9042_o & n9020_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9048_o = challenge == 8'b10101111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9049_o = sortie_ro[175];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9050_o = n9061_o ? n9049_o : n9032_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9052_o = n9063_o ? 1'b1 : n9034_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9056_o = n9064_o ? 1'b0 : n9038_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9057_o = n9038_o & n9048_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9059_o = n9038_o & n9048_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9060_o = n9038_o & n9048_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9061_o = n9057_o & n9038_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9063_o = n9059_o & n9038_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9064_o = n9060_o & n9038_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9066_o = challenge == 8'b10110000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9067_o = sortie_ro[176];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9068_o = n9079_o ? n9067_o : n9050_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9070_o = n9081_o ? 1'b1 : n9052_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9074_o = n9082_o ? 1'b0 : n9056_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9075_o = n9056_o & n9066_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9077_o = n9056_o & n9066_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9078_o = n9056_o & n9066_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9079_o = n9075_o & n9056_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9081_o = n9077_o & n9056_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9082_o = n9078_o & n9056_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9084_o = challenge == 8'b10110001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9085_o = sortie_ro[177];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9086_o = n9097_o ? n9085_o : n9068_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9088_o = n9099_o ? 1'b1 : n9070_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9092_o = n9100_o ? 1'b0 : n9074_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9093_o = n9074_o & n9084_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9095_o = n9074_o & n9084_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9096_o = n9074_o & n9084_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9097_o = n9093_o & n9074_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9099_o = n9095_o & n9074_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9100_o = n9096_o & n9074_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9102_o = challenge == 8'b10110010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9103_o = sortie_ro[178];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9104_o = n9115_o ? n9103_o : n9086_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9106_o = n9117_o ? 1'b1 : n9088_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9110_o = n9118_o ? 1'b0 : n9092_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9111_o = n9092_o & n9102_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9113_o = n9092_o & n9102_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9114_o = n9092_o & n9102_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9115_o = n9111_o & n9092_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9117_o = n9113_o & n9092_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9118_o = n9114_o & n9092_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9120_o = challenge == 8'b10110011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9121_o = sortie_ro[179];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9122_o = n9133_o ? n9121_o : n9104_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9124_o = n9135_o ? 1'b1 : n9106_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9128_o = n9136_o ? 1'b0 : n9110_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9129_o = n9110_o & n9120_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9131_o = n9110_o & n9120_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9132_o = n9110_o & n9120_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9133_o = n9129_o & n9110_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9135_o = n9131_o & n9110_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9136_o = n9132_o & n9110_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9138_o = challenge == 8'b10110100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9139_o = sortie_ro[180];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9140_o = n9151_o ? n9139_o : n9122_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9142_o = n9153_o ? 1'b1 : n9124_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9146_o = n9154_o ? 1'b0 : n9128_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9147_o = n9128_o & n9138_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9149_o = n9128_o & n9138_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9150_o = n9128_o & n9138_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9151_o = n9147_o & n9128_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9153_o = n9149_o & n9128_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9154_o = n9150_o & n9128_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9156_o = challenge == 8'b10110101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9157_o = sortie_ro[181];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9158_o = n9169_o ? n9157_o : n9140_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9160_o = n9171_o ? 1'b1 : n9142_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9164_o = n9172_o ? 1'b0 : n9146_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9165_o = n9146_o & n9156_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9167_o = n9146_o & n9156_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9168_o = n9146_o & n9156_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9169_o = n9165_o & n9146_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9171_o = n9167_o & n9146_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9172_o = n9168_o & n9146_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9174_o = challenge == 8'b10110110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9175_o = sortie_ro[182];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9176_o = n9187_o ? n9175_o : n9158_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9178_o = n9189_o ? 1'b1 : n9160_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9182_o = n9190_o ? 1'b0 : n9164_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9183_o = n9164_o & n9174_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9185_o = n9164_o & n9174_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9186_o = n9164_o & n9174_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9187_o = n9183_o & n9164_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9189_o = n9185_o & n9164_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9190_o = n9186_o & n9164_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9192_o = challenge == 8'b10110111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9193_o = sortie_ro[183];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9194_o = n9205_o ? n9193_o : n9176_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9196_o = n9207_o ? 1'b1 : n9178_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9200_o = n9208_o ? 1'b0 : n9182_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9201_o = n9182_o & n9192_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9203_o = n9182_o & n9192_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9204_o = n9182_o & n9192_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9205_o = n9201_o & n9182_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9207_o = n9203_o & n9182_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9208_o = n9204_o & n9182_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9210_o = challenge == 8'b10111000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9211_o = sortie_ro[184];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9212_o = n9223_o ? n9211_o : n9194_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9214_o = n9225_o ? 1'b1 : n9196_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9218_o = n9226_o ? 1'b0 : n9200_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9219_o = n9200_o & n9210_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9221_o = n9200_o & n9210_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9222_o = n9200_o & n9210_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9223_o = n9219_o & n9200_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9225_o = n9221_o & n9200_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9226_o = n9222_o & n9200_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9228_o = challenge == 8'b10111001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9229_o = sortie_ro[185];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9230_o = n9241_o ? n9229_o : n9212_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9232_o = n9243_o ? 1'b1 : n9214_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9236_o = n9244_o ? 1'b0 : n9218_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9237_o = n9218_o & n9228_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9239_o = n9218_o & n9228_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9240_o = n9218_o & n9228_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9241_o = n9237_o & n9218_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9243_o = n9239_o & n9218_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9244_o = n9240_o & n9218_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9246_o = challenge == 8'b10111010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9247_o = sortie_ro[186];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9248_o = n9259_o ? n9247_o : n9230_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9250_o = n9261_o ? 1'b1 : n9232_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9254_o = n9262_o ? 1'b0 : n9236_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9255_o = n9236_o & n9246_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9257_o = n9236_o & n9246_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9258_o = n9236_o & n9246_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9259_o = n9255_o & n9236_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9261_o = n9257_o & n9236_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9262_o = n9258_o & n9236_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9264_o = challenge == 8'b10111011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9265_o = sortie_ro[187];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9266_o = n9277_o ? n9265_o : n9248_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9268_o = n9279_o ? 1'b1 : n9250_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9272_o = n9280_o ? 1'b0 : n9254_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9273_o = n9254_o & n9264_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9275_o = n9254_o & n9264_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9276_o = n9254_o & n9264_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9277_o = n9273_o & n9254_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9279_o = n9275_o & n9254_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9280_o = n9276_o & n9254_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9282_o = challenge == 8'b10111100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9283_o = sortie_ro[188];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9284_o = n9295_o ? n9283_o : n9266_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9286_o = n9297_o ? 1'b1 : n9268_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9290_o = n9298_o ? 1'b0 : n9272_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9291_o = n9272_o & n9282_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9293_o = n9272_o & n9282_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9294_o = n9272_o & n9282_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9295_o = n9291_o & n9272_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9297_o = n9293_o & n9272_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9298_o = n9294_o & n9272_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9300_o = challenge == 8'b10111101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9301_o = sortie_ro[189];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9302_o = n9313_o ? n9301_o : n9284_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9304_o = n9315_o ? 1'b1 : n9286_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9308_o = n9316_o ? 1'b0 : n9290_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9309_o = n9290_o & n9300_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9311_o = n9290_o & n9300_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9312_o = n9290_o & n9300_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9313_o = n9309_o & n9290_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9315_o = n9311_o & n9290_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9316_o = n9312_o & n9290_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9318_o = challenge == 8'b10111110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9319_o = sortie_ro[190];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9320_o = n9331_o ? n9319_o : n9302_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9322_o = n9333_o ? 1'b1 : n9304_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9326_o = n9334_o ? 1'b0 : n9308_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9327_o = n9308_o & n9318_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9329_o = n9308_o & n9318_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9330_o = n9308_o & n9318_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9331_o = n9327_o & n9308_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9333_o = n9329_o & n9308_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9334_o = n9330_o & n9308_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9336_o = challenge == 8'b10111111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9337_o = sortie_ro[191];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9338_o = n9349_o ? n9337_o : n9320_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9340_o = n9351_o ? 1'b1 : n9322_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9344_o = n9352_o ? 1'b0 : n9326_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9345_o = n9326_o & n9336_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9347_o = n9326_o & n9336_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9348_o = n9326_o & n9336_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9349_o = n9345_o & n9326_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9351_o = n9347_o & n9326_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9352_o = n9348_o & n9326_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9354_o = challenge == 8'b11000000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9355_o = sortie_ro[192];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9356_o = n9367_o ? n9355_o : n9338_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9358_o = n9369_o ? 1'b1 : n9340_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9362_o = n9370_o ? 1'b0 : n9344_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9363_o = n9344_o & n9354_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9365_o = n9344_o & n9354_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9366_o = n9344_o & n9354_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9367_o = n9363_o & n9344_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9369_o = n9365_o & n9344_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9370_o = n9366_o & n9344_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9372_o = challenge == 8'b11000001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9373_o = sortie_ro[193];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9374_o = n9385_o ? n9373_o : n9356_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9376_o = n9387_o ? 1'b1 : n9358_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9380_o = n9388_o ? 1'b0 : n9362_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9381_o = n9362_o & n9372_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9383_o = n9362_o & n9372_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9384_o = n9362_o & n9372_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9385_o = n9381_o & n9362_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9387_o = n9383_o & n9362_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9388_o = n9384_o & n9362_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9390_o = challenge == 8'b11000010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9391_o = sortie_ro[194];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9392_o = n9403_o ? n9391_o : n9374_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9394_o = n9405_o ? 1'b1 : n9376_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9398_o = n9406_o ? 1'b0 : n9380_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9399_o = n9380_o & n9390_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9401_o = n9380_o & n9390_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9402_o = n9380_o & n9390_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9403_o = n9399_o & n9380_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9405_o = n9401_o & n9380_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9406_o = n9402_o & n9380_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9408_o = challenge == 8'b11000011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9409_o = sortie_ro[195];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9410_o = n9421_o ? n9409_o : n9392_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9412_o = n9423_o ? 1'b1 : n9394_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9416_o = n9424_o ? 1'b0 : n9398_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9417_o = n9398_o & n9408_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9419_o = n9398_o & n9408_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9420_o = n9398_o & n9408_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9421_o = n9417_o & n9398_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9423_o = n9419_o & n9398_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9424_o = n9420_o & n9398_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9426_o = challenge == 8'b11000100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9427_o = sortie_ro[196];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9428_o = n9439_o ? n9427_o : n9410_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9430_o = n9441_o ? 1'b1 : n9412_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9434_o = n9442_o ? 1'b0 : n9416_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9435_o = n9416_o & n9426_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9437_o = n9416_o & n9426_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9438_o = n9416_o & n9426_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9439_o = n9435_o & n9416_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9441_o = n9437_o & n9416_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9442_o = n9438_o & n9416_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9444_o = challenge == 8'b11000101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9445_o = sortie_ro[197];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9446_o = n9457_o ? n9445_o : n9428_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9448_o = n9459_o ? 1'b1 : n9430_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9452_o = n9460_o ? 1'b0 : n9434_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9453_o = n9434_o & n9444_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9455_o = n9434_o & n9444_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9456_o = n9434_o & n9444_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9457_o = n9453_o & n9434_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9459_o = n9455_o & n9434_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9460_o = n9456_o & n9434_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9462_o = challenge == 8'b11000110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9463_o = sortie_ro[198];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9464_o = n9475_o ? n9463_o : n9446_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9466_o = n9477_o ? 1'b1 : n9448_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9470_o = n9478_o ? 1'b0 : n9452_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9471_o = n9452_o & n9462_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9473_o = n9452_o & n9462_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9474_o = n9452_o & n9462_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9475_o = n9471_o & n9452_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9477_o = n9473_o & n9452_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9478_o = n9474_o & n9452_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9480_o = challenge == 8'b11000111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9481_o = sortie_ro[199];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9482_o = n9493_o ? n9481_o : n9464_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9484_o = n9495_o ? 1'b1 : n9466_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9488_o = n9496_o ? 1'b0 : n9470_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9489_o = n9470_o & n9480_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9491_o = n9470_o & n9480_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9492_o = n9470_o & n9480_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9493_o = n9489_o & n9470_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9495_o = n9491_o & n9470_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9496_o = n9492_o & n9470_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9498_o = challenge == 8'b11001000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9499_o = sortie_ro[200];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9500_o = n9511_o ? n9499_o : n9482_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9502_o = n9513_o ? 1'b1 : n9484_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9506_o = n9514_o ? 1'b0 : n9488_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9507_o = n9488_o & n9498_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9509_o = n9488_o & n9498_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9510_o = n9488_o & n9498_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9511_o = n9507_o & n9488_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9513_o = n9509_o & n9488_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9514_o = n9510_o & n9488_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9516_o = challenge == 8'b11001001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9517_o = sortie_ro[201];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9518_o = n9529_o ? n9517_o : n9500_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9520_o = n9531_o ? 1'b1 : n9502_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9524_o = n9532_o ? 1'b0 : n9506_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9525_o = n9506_o & n9516_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9527_o = n9506_o & n9516_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9528_o = n9506_o & n9516_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9529_o = n9525_o & n9506_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9531_o = n9527_o & n9506_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9532_o = n9528_o & n9506_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9534_o = challenge == 8'b11001010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9535_o = sortie_ro[202];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9536_o = n9547_o ? n9535_o : n9518_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9538_o = n9549_o ? 1'b1 : n9520_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9542_o = n9550_o ? 1'b0 : n9524_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9543_o = n9524_o & n9534_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9545_o = n9524_o & n9534_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9546_o = n9524_o & n9534_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9547_o = n9543_o & n9524_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9549_o = n9545_o & n9524_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9550_o = n9546_o & n9524_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9552_o = challenge == 8'b11001011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9553_o = sortie_ro[203];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9554_o = n9565_o ? n9553_o : n9536_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9556_o = n9567_o ? 1'b1 : n9538_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9560_o = n9568_o ? 1'b0 : n9542_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9561_o = n9542_o & n9552_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9563_o = n9542_o & n9552_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9564_o = n9542_o & n9552_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9565_o = n9561_o & n9542_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9567_o = n9563_o & n9542_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9568_o = n9564_o & n9542_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9570_o = challenge == 8'b11001100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9571_o = sortie_ro[204];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9572_o = n9583_o ? n9571_o : n9554_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9574_o = n9585_o ? 1'b1 : n9556_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9578_o = n9586_o ? 1'b0 : n9560_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9579_o = n9560_o & n9570_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9581_o = n9560_o & n9570_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9582_o = n9560_o & n9570_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9583_o = n9579_o & n9560_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9585_o = n9581_o & n9560_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9586_o = n9582_o & n9560_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9588_o = challenge == 8'b11001101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9589_o = sortie_ro[205];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9590_o = n9601_o ? n9589_o : n9572_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9592_o = n9603_o ? 1'b1 : n9574_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9596_o = n9604_o ? 1'b0 : n9578_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9597_o = n9578_o & n9588_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9599_o = n9578_o & n9588_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9600_o = n9578_o & n9588_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9601_o = n9597_o & n9578_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9603_o = n9599_o & n9578_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9604_o = n9600_o & n9578_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9606_o = challenge == 8'b11001110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9607_o = sortie_ro[206];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9608_o = n9619_o ? n9607_o : n9590_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9610_o = n9621_o ? 1'b1 : n9592_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9614_o = n9622_o ? 1'b0 : n9596_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9615_o = n9596_o & n9606_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9617_o = n9596_o & n9606_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9618_o = n9596_o & n9606_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9619_o = n9615_o & n9596_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9621_o = n9617_o & n9596_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9622_o = n9618_o & n9596_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9624_o = challenge == 8'b11001111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9625_o = sortie_ro[207];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9626_o = n9637_o ? n9625_o : n9608_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9628_o = n9639_o ? 1'b1 : n9610_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9632_o = n9640_o ? 1'b0 : n9614_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9633_o = n9614_o & n9624_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9635_o = n9614_o & n9624_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9636_o = n9614_o & n9624_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9637_o = n9633_o & n9614_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9639_o = n9635_o & n9614_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9640_o = n9636_o & n9614_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9642_o = challenge == 8'b11010000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9643_o = sortie_ro[208];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9644_o = n9655_o ? n9643_o : n9626_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9646_o = n9657_o ? 1'b1 : n9628_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9650_o = n9658_o ? 1'b0 : n9632_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9651_o = n9632_o & n9642_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9653_o = n9632_o & n9642_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9654_o = n9632_o & n9642_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9655_o = n9651_o & n9632_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9657_o = n9653_o & n9632_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9658_o = n9654_o & n9632_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9660_o = challenge == 8'b11010001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9661_o = sortie_ro[209];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9662_o = n9673_o ? n9661_o : n9644_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9664_o = n9675_o ? 1'b1 : n9646_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9668_o = n9676_o ? 1'b0 : n9650_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9669_o = n9650_o & n9660_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9671_o = n9650_o & n9660_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9672_o = n9650_o & n9660_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9673_o = n9669_o & n9650_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9675_o = n9671_o & n9650_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9676_o = n9672_o & n9650_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9678_o = challenge == 8'b11010010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9679_o = sortie_ro[210];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9680_o = n9691_o ? n9679_o : n9662_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9682_o = n9693_o ? 1'b1 : n9664_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9686_o = n9694_o ? 1'b0 : n9668_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9687_o = n9668_o & n9678_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9689_o = n9668_o & n9678_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9690_o = n9668_o & n9678_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9691_o = n9687_o & n9668_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9693_o = n9689_o & n9668_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9694_o = n9690_o & n9668_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9696_o = challenge == 8'b11010011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9697_o = sortie_ro[211];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9698_o = n9709_o ? n9697_o : n9680_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9700_o = n9711_o ? 1'b1 : n9682_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9704_o = n9712_o ? 1'b0 : n9686_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9705_o = n9686_o & n9696_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9707_o = n9686_o & n9696_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9708_o = n9686_o & n9696_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9709_o = n9705_o & n9686_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9711_o = n9707_o & n9686_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9712_o = n9708_o & n9686_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9714_o = challenge == 8'b11010100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9715_o = sortie_ro[212];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9716_o = n9727_o ? n9715_o : n9698_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9718_o = n9729_o ? 1'b1 : n9700_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9722_o = n9730_o ? 1'b0 : n9704_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9723_o = n9704_o & n9714_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9725_o = n9704_o & n9714_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9726_o = n9704_o & n9714_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9727_o = n9723_o & n9704_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9729_o = n9725_o & n9704_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9730_o = n9726_o & n9704_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9732_o = challenge == 8'b11010101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9733_o = sortie_ro[213];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9734_o = n9745_o ? n9733_o : n9716_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9736_o = n9747_o ? 1'b1 : n9718_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9740_o = n9748_o ? 1'b0 : n9722_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9741_o = n9722_o & n9732_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9743_o = n9722_o & n9732_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9744_o = n9722_o & n9732_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9745_o = n9741_o & n9722_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9747_o = n9743_o & n9722_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9748_o = n9744_o & n9722_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9750_o = challenge == 8'b11010110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9751_o = sortie_ro[214];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9752_o = n9763_o ? n9751_o : n9734_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9754_o = n9765_o ? 1'b1 : n9736_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9758_o = n9766_o ? 1'b0 : n9740_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9759_o = n9740_o & n9750_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9761_o = n9740_o & n9750_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9762_o = n9740_o & n9750_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9763_o = n9759_o & n9740_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9765_o = n9761_o & n9740_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9766_o = n9762_o & n9740_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9768_o = challenge == 8'b11010111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9769_o = sortie_ro[215];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9770_o = n9781_o ? n9769_o : n9752_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9772_o = n9783_o ? 1'b1 : n9754_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9776_o = n9784_o ? 1'b0 : n9758_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9777_o = n9758_o & n9768_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9779_o = n9758_o & n9768_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9780_o = n9758_o & n9768_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9781_o = n9777_o & n9758_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9783_o = n9779_o & n9758_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9784_o = n9780_o & n9758_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9786_o = challenge == 8'b11011000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9787_o = sortie_ro[216];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9788_o = n9799_o ? n9787_o : n9770_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9790_o = n9801_o ? 1'b1 : n9772_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9794_o = n9802_o ? 1'b0 : n9776_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9795_o = n9776_o & n9786_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9797_o = n9776_o & n9786_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9798_o = n9776_o & n9786_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9799_o = n9795_o & n9776_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9801_o = n9797_o & n9776_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9802_o = n9798_o & n9776_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9804_o = challenge == 8'b11011001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9805_o = sortie_ro[217];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9806_o = n9817_o ? n9805_o : n9788_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9808_o = n9819_o ? 1'b1 : n9790_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9812_o = n9820_o ? 1'b0 : n9794_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9813_o = n9794_o & n9804_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9815_o = n9794_o & n9804_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9816_o = n9794_o & n9804_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9817_o = n9813_o & n9794_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9819_o = n9815_o & n9794_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9820_o = n9816_o & n9794_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9822_o = challenge == 8'b11011010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9823_o = sortie_ro[218];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9824_o = n9835_o ? n9823_o : n9806_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9826_o = n9837_o ? 1'b1 : n9808_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9830_o = n9838_o ? 1'b0 : n9812_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9831_o = n9812_o & n9822_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9833_o = n9812_o & n9822_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9834_o = n9812_o & n9822_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9835_o = n9831_o & n9812_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9837_o = n9833_o & n9812_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9838_o = n9834_o & n9812_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9840_o = challenge == 8'b11011011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9841_o = sortie_ro[219];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9842_o = n9853_o ? n9841_o : n9824_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9844_o = n9855_o ? 1'b1 : n9826_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9848_o = n9856_o ? 1'b0 : n9830_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9849_o = n9830_o & n9840_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9851_o = n9830_o & n9840_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9852_o = n9830_o & n9840_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9853_o = n9849_o & n9830_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9855_o = n9851_o & n9830_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9856_o = n9852_o & n9830_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9858_o = challenge == 8'b11011100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9859_o = sortie_ro[220];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9860_o = n9871_o ? n9859_o : n9842_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9862_o = n9873_o ? 1'b1 : n9844_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9866_o = n9874_o ? 1'b0 : n9848_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9867_o = n9848_o & n9858_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9869_o = n9848_o & n9858_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9870_o = n9848_o & n9858_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9871_o = n9867_o & n9848_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9873_o = n9869_o & n9848_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9874_o = n9870_o & n9848_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9876_o = challenge == 8'b11011101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9877_o = sortie_ro[221];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9878_o = n9889_o ? n9877_o : n9860_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9880_o = n9891_o ? 1'b1 : n9862_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9884_o = n9892_o ? 1'b0 : n9866_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9885_o = n9866_o & n9876_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9887_o = n9866_o & n9876_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9888_o = n9866_o & n9876_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9889_o = n9885_o & n9866_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9891_o = n9887_o & n9866_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9892_o = n9888_o & n9866_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9894_o = challenge == 8'b11011110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9895_o = sortie_ro[222];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9896_o = n9907_o ? n9895_o : n9878_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9898_o = n9909_o ? 1'b1 : n9880_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9902_o = n9910_o ? 1'b0 : n9884_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9903_o = n9884_o & n9894_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9905_o = n9884_o & n9894_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9906_o = n9884_o & n9894_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9907_o = n9903_o & n9884_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9909_o = n9905_o & n9884_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9910_o = n9906_o & n9884_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9912_o = challenge == 8'b11011111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9913_o = sortie_ro[223];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9914_o = n9925_o ? n9913_o : n9896_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9916_o = n9927_o ? 1'b1 : n9898_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9920_o = n9928_o ? 1'b0 : n9902_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9921_o = n9902_o & n9912_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9923_o = n9902_o & n9912_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9924_o = n9902_o & n9912_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9925_o = n9921_o & n9902_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9927_o = n9923_o & n9902_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9928_o = n9924_o & n9902_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9930_o = challenge == 8'b11100000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9931_o = sortie_ro[224];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9932_o = n9943_o ? n9931_o : n9914_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9934_o = n9945_o ? 1'b1 : n9916_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9938_o = n9946_o ? 1'b0 : n9920_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9939_o = n9920_o & n9930_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9941_o = n9920_o & n9930_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9942_o = n9920_o & n9930_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9943_o = n9939_o & n9920_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9945_o = n9941_o & n9920_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9946_o = n9942_o & n9920_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9948_o = challenge == 8'b11100001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9949_o = sortie_ro[225];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9950_o = n9961_o ? n9949_o : n9932_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9952_o = n9963_o ? 1'b1 : n9934_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9956_o = n9964_o ? 1'b0 : n9938_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9957_o = n9938_o & n9948_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9959_o = n9938_o & n9948_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9960_o = n9938_o & n9948_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9961_o = n9957_o & n9938_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9963_o = n9959_o & n9938_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9964_o = n9960_o & n9938_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9966_o = challenge == 8'b11100010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9967_o = sortie_ro[226];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9968_o = n9979_o ? n9967_o : n9950_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9970_o = n9981_o ? 1'b1 : n9952_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9974_o = n9982_o ? 1'b0 : n9956_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9975_o = n9956_o & n9966_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9977_o = n9956_o & n9966_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9978_o = n9956_o & n9966_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9979_o = n9975_o & n9956_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9981_o = n9977_o & n9956_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9982_o = n9978_o & n9956_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n9984_o = challenge == 8'b11100011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n9985_o = sortie_ro[227];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9986_o = n9997_o ? n9985_o : n9968_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9988_o = n9999_o ? 1'b1 : n9970_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9992_o = n10000_o ? 1'b0 : n9974_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9993_o = n9974_o & n9984_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9995_o = n9974_o & n9984_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9996_o = n9974_o & n9984_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9997_o = n9993_o & n9974_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n9999_o = n9995_o & n9974_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10000_o = n9996_o & n9974_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10002_o = challenge == 8'b11100100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10003_o = sortie_ro[228];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10004_o = n10015_o ? n10003_o : n9986_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10006_o = n10017_o ? 1'b1 : n9988_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10010_o = n10018_o ? 1'b0 : n9992_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10011_o = n9992_o & n10002_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10013_o = n9992_o & n10002_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10014_o = n9992_o & n10002_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10015_o = n10011_o & n9992_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10017_o = n10013_o & n9992_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10018_o = n10014_o & n9992_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10020_o = challenge == 8'b11100101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10021_o = sortie_ro[229];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10022_o = n10033_o ? n10021_o : n10004_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10024_o = n10035_o ? 1'b1 : n10006_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10028_o = n10036_o ? 1'b0 : n10010_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10029_o = n10010_o & n10020_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10031_o = n10010_o & n10020_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10032_o = n10010_o & n10020_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10033_o = n10029_o & n10010_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10035_o = n10031_o & n10010_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10036_o = n10032_o & n10010_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10038_o = challenge == 8'b11100110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10039_o = sortie_ro[230];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10040_o = n10051_o ? n10039_o : n10022_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10042_o = n10053_o ? 1'b1 : n10024_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10046_o = n10054_o ? 1'b0 : n10028_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10047_o = n10028_o & n10038_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10049_o = n10028_o & n10038_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10050_o = n10028_o & n10038_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10051_o = n10047_o & n10028_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10053_o = n10049_o & n10028_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10054_o = n10050_o & n10028_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10056_o = challenge == 8'b11100111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10057_o = sortie_ro[231];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10058_o = n10069_o ? n10057_o : n10040_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10060_o = n10071_o ? 1'b1 : n10042_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10064_o = n10072_o ? 1'b0 : n10046_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10065_o = n10046_o & n10056_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10067_o = n10046_o & n10056_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10068_o = n10046_o & n10056_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10069_o = n10065_o & n10046_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10071_o = n10067_o & n10046_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10072_o = n10068_o & n10046_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10074_o = challenge == 8'b11101000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10075_o = sortie_ro[232];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10076_o = n10087_o ? n10075_o : n10058_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10078_o = n10089_o ? 1'b1 : n10060_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10082_o = n10090_o ? 1'b0 : n10064_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10083_o = n10064_o & n10074_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10085_o = n10064_o & n10074_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10086_o = n10064_o & n10074_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10087_o = n10083_o & n10064_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10089_o = n10085_o & n10064_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10090_o = n10086_o & n10064_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10092_o = challenge == 8'b11101001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10093_o = sortie_ro[233];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10094_o = n10105_o ? n10093_o : n10076_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10096_o = n10107_o ? 1'b1 : n10078_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10100_o = n10108_o ? 1'b0 : n10082_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10101_o = n10082_o & n10092_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10103_o = n10082_o & n10092_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10104_o = n10082_o & n10092_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10105_o = n10101_o & n10082_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10107_o = n10103_o & n10082_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10108_o = n10104_o & n10082_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10110_o = challenge == 8'b11101010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10111_o = sortie_ro[234];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10112_o = n10123_o ? n10111_o : n10094_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10114_o = n10125_o ? 1'b1 : n10096_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10118_o = n10126_o ? 1'b0 : n10100_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10119_o = n10100_o & n10110_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10121_o = n10100_o & n10110_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10122_o = n10100_o & n10110_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10123_o = n10119_o & n10100_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10125_o = n10121_o & n10100_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10126_o = n10122_o & n10100_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10128_o = challenge == 8'b11101011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10129_o = sortie_ro[235];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10130_o = n10141_o ? n10129_o : n10112_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10132_o = n10143_o ? 1'b1 : n10114_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10136_o = n10144_o ? 1'b0 : n10118_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10137_o = n10118_o & n10128_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10139_o = n10118_o & n10128_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10140_o = n10118_o & n10128_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10141_o = n10137_o & n10118_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10143_o = n10139_o & n10118_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10144_o = n10140_o & n10118_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10146_o = challenge == 8'b11101100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10147_o = sortie_ro[236];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10148_o = n10159_o ? n10147_o : n10130_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10150_o = n10161_o ? 1'b1 : n10132_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10154_o = n10162_o ? 1'b0 : n10136_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10155_o = n10136_o & n10146_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10157_o = n10136_o & n10146_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10158_o = n10136_o & n10146_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10159_o = n10155_o & n10136_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10161_o = n10157_o & n10136_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10162_o = n10158_o & n10136_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10164_o = challenge == 8'b11101101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10165_o = sortie_ro[237];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10166_o = n10177_o ? n10165_o : n10148_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10168_o = n10179_o ? 1'b1 : n10150_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10172_o = n10180_o ? 1'b0 : n10154_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10173_o = n10154_o & n10164_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10175_o = n10154_o & n10164_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10176_o = n10154_o & n10164_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10177_o = n10173_o & n10154_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10179_o = n10175_o & n10154_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10180_o = n10176_o & n10154_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10182_o = challenge == 8'b11101110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10183_o = sortie_ro[238];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10184_o = n10195_o ? n10183_o : n10166_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10186_o = n10197_o ? 1'b1 : n10168_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10190_o = n10198_o ? 1'b0 : n10172_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10191_o = n10172_o & n10182_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10193_o = n10172_o & n10182_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10194_o = n10172_o & n10182_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10195_o = n10191_o & n10172_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10197_o = n10193_o & n10172_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10198_o = n10194_o & n10172_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10200_o = challenge == 8'b11101111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10201_o = sortie_ro[239];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10202_o = n10213_o ? n10201_o : n10184_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10204_o = n10215_o ? 1'b1 : n10186_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10208_o = n10216_o ? 1'b0 : n10190_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10209_o = n10190_o & n10200_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10211_o = n10190_o & n10200_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10212_o = n10190_o & n10200_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10213_o = n10209_o & n10190_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10215_o = n10211_o & n10190_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10216_o = n10212_o & n10190_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10218_o = challenge == 8'b11110000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10219_o = sortie_ro[240];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10220_o = n10231_o ? n10219_o : n10202_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10222_o = n10233_o ? 1'b1 : n10204_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10226_o = n10234_o ? 1'b0 : n10208_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10227_o = n10208_o & n10218_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10229_o = n10208_o & n10218_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10230_o = n10208_o & n10218_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10231_o = n10227_o & n10208_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10233_o = n10229_o & n10208_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10234_o = n10230_o & n10208_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10236_o = challenge == 8'b11110001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10237_o = sortie_ro[241];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10238_o = n10249_o ? n10237_o : n10220_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10240_o = n10251_o ? 1'b1 : n10222_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10244_o = n10252_o ? 1'b0 : n10226_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10245_o = n10226_o & n10236_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10247_o = n10226_o & n10236_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10248_o = n10226_o & n10236_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10249_o = n10245_o & n10226_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10251_o = n10247_o & n10226_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10252_o = n10248_o & n10226_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10254_o = challenge == 8'b11110010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10255_o = sortie_ro[242];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10256_o = n10267_o ? n10255_o : n10238_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10258_o = n10269_o ? 1'b1 : n10240_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10262_o = n10270_o ? 1'b0 : n10244_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10263_o = n10244_o & n10254_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10265_o = n10244_o & n10254_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10266_o = n10244_o & n10254_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10267_o = n10263_o & n10244_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10269_o = n10265_o & n10244_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10270_o = n10266_o & n10244_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10272_o = challenge == 8'b11110011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10273_o = sortie_ro[243];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10274_o = n10285_o ? n10273_o : n10256_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10276_o = n10287_o ? 1'b1 : n10258_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10280_o = n10288_o ? 1'b0 : n10262_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10281_o = n10262_o & n10272_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10283_o = n10262_o & n10272_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10284_o = n10262_o & n10272_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10285_o = n10281_o & n10262_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10287_o = n10283_o & n10262_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10288_o = n10284_o & n10262_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10290_o = challenge == 8'b11110100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10291_o = sortie_ro[244];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10292_o = n10303_o ? n10291_o : n10274_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10294_o = n10305_o ? 1'b1 : n10276_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10298_o = n10306_o ? 1'b0 : n10280_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10299_o = n10280_o & n10290_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10301_o = n10280_o & n10290_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10302_o = n10280_o & n10290_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10303_o = n10299_o & n10280_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10305_o = n10301_o & n10280_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10306_o = n10302_o & n10280_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10308_o = challenge == 8'b11110101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10309_o = sortie_ro[245];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10310_o = n10321_o ? n10309_o : n10292_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10312_o = n10323_o ? 1'b1 : n10294_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10316_o = n10324_o ? 1'b0 : n10298_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10317_o = n10298_o & n10308_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10319_o = n10298_o & n10308_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10320_o = n10298_o & n10308_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10321_o = n10317_o & n10298_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10323_o = n10319_o & n10298_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10324_o = n10320_o & n10298_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10326_o = challenge == 8'b11110110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10327_o = sortie_ro[246];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10328_o = n10339_o ? n10327_o : n10310_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10330_o = n10341_o ? 1'b1 : n10312_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10334_o = n10342_o ? 1'b0 : n10316_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10335_o = n10316_o & n10326_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10337_o = n10316_o & n10326_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10338_o = n10316_o & n10326_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10339_o = n10335_o & n10316_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10341_o = n10337_o & n10316_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10342_o = n10338_o & n10316_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10344_o = challenge == 8'b11110111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10345_o = sortie_ro[247];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10346_o = n10357_o ? n10345_o : n10328_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10348_o = n10359_o ? 1'b1 : n10330_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10352_o = n10360_o ? 1'b0 : n10334_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10353_o = n10334_o & n10344_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10355_o = n10334_o & n10344_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10356_o = n10334_o & n10344_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10357_o = n10353_o & n10334_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10359_o = n10355_o & n10334_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10360_o = n10356_o & n10334_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10362_o = challenge == 8'b11111000;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10363_o = sortie_ro[248];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10364_o = n10375_o ? n10363_o : n10346_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10366_o = n10377_o ? 1'b1 : n10348_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10370_o = n10378_o ? 1'b0 : n10352_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10371_o = n10352_o & n10362_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10373_o = n10352_o & n10362_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10374_o = n10352_o & n10362_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10375_o = n10371_o & n10352_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10377_o = n10373_o & n10352_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10378_o = n10374_o & n10352_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10380_o = challenge == 8'b11111001;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10381_o = sortie_ro[249];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10382_o = n10393_o ? n10381_o : n10364_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10384_o = n10395_o ? 1'b1 : n10366_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10388_o = n10396_o ? 1'b0 : n10370_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10389_o = n10370_o & n10380_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10391_o = n10370_o & n10380_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10392_o = n10370_o & n10380_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10393_o = n10389_o & n10370_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10395_o = n10391_o & n10370_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10396_o = n10392_o & n10370_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10398_o = challenge == 8'b11111010;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10399_o = sortie_ro[250];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10400_o = n10411_o ? n10399_o : n10382_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10402_o = n10413_o ? 1'b1 : n10384_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10406_o = n10414_o ? 1'b0 : n10388_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10407_o = n10388_o & n10398_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10409_o = n10388_o & n10398_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10410_o = n10388_o & n10398_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10411_o = n10407_o & n10388_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10413_o = n10409_o & n10388_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10414_o = n10410_o & n10388_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10416_o = challenge == 8'b11111011;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10417_o = sortie_ro[251];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10418_o = n10429_o ? n10417_o : n10400_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10420_o = n10431_o ? 1'b1 : n10402_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10424_o = n10432_o ? 1'b0 : n10406_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10425_o = n10406_o & n10416_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10427_o = n10406_o & n10416_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10428_o = n10406_o & n10416_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10429_o = n10425_o & n10406_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10431_o = n10427_o & n10406_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10432_o = n10428_o & n10406_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10434_o = challenge == 8'b11111100;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10435_o = sortie_ro[252];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10436_o = n10447_o ? n10435_o : n10418_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10438_o = n10449_o ? 1'b1 : n10420_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10442_o = n10450_o ? 1'b0 : n10424_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10443_o = n10424_o & n10434_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10445_o = n10424_o & n10434_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10446_o = n10424_o & n10434_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10447_o = n10443_o & n10424_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10449_o = n10445_o & n10424_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10450_o = n10446_o & n10424_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10452_o = challenge == 8'b11111101;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10453_o = sortie_ro[253];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10454_o = n10465_o ? n10453_o : n10436_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10456_o = n10467_o ? 1'b1 : n10438_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10460_o = n10468_o ? 1'b0 : n10442_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10461_o = n10442_o & n10452_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10463_o = n10442_o & n10452_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10464_o = n10442_o & n10452_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10465_o = n10461_o & n10442_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10467_o = n10463_o & n10442_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10468_o = n10464_o & n10442_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10470_o = challenge == 8'b11111110;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10471_o = sortie_ro[254];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10472_o = n10483_o ? n10471_o : n10454_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10474_o = n10485_o ? 1'b1 : n10456_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10478_o = n10486_o ? 1'b0 : n10460_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10479_o = n10460_o & n10470_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10481_o = n10460_o & n10470_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10482_o = n10460_o & n10470_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10483_o = n10479_o & n10460_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10485_o = n10481_o & n10460_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10486_o = n10482_o & n10460_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:22  */
  assign n10488_o = challenge == 8'b11111111;
  /* RTL_PUF/vhdl/ro_array.vhd:49:32  */
  assign n10489_o = sortie_ro[255];
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10490_o = n10501_o ? n10489_o : n10472_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10492_o = n10503_o ? 1'b1 : n10474_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10497_o = n10478_o & n10488_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10499_o = n10478_o & n10488_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10501_o = n10497_o & n10478_o;
  /* RTL_PUF/vhdl/ro_array.vhd:48:9  */
  assign n10503_o = n10499_o & n10478_o;
  /* RTL_PUF/vhdl/ro_array.vhd:54:8  */
  assign n10505_o = ~n10492_o;
  /* RTL_PUF/vhdl/ro_array.vhd:54:5  */
  assign n10507_o = n10505_o ? 1'b0 : n10490_o;
  assign n10765_o = {inverseur_n256_ringoscillator_n5894, inverseur_n255_ringoscillator_n5890, inverseur_n254_ringoscillator_n5886, inverseur_n253_ringoscillator_n5882, inverseur_n252_ringoscillator_n5878, inverseur_n251_ringoscillator_n5874, inverseur_n250_ringoscillator_n5870, inverseur_n249_ringoscillator_n5866, inverseur_n248_ringoscillator_n5862, inverseur_n247_ringoscillator_n5858, inverseur_n246_ringoscillator_n5854, inverseur_n245_ringoscillator_n5850, inverseur_n244_ringoscillator_n5846, inverseur_n243_ringoscillator_n5842, inverseur_n242_ringoscillator_n5838, inverseur_n241_ringoscillator_n5834, inverseur_n240_ringoscillator_n5830, inverseur_n239_ringoscillator_n5826, inverseur_n238_ringoscillator_n5822, inverseur_n237_ringoscillator_n5818, inverseur_n236_ringoscillator_n5814, inverseur_n235_ringoscillator_n5810, inverseur_n234_ringoscillator_n5806, inverseur_n233_ringoscillator_n5802, inverseur_n232_ringoscillator_n5798, inverseur_n231_ringoscillator_n5794, inverseur_n230_ringoscillator_n5790, inverseur_n229_ringoscillator_n5786, inverseur_n228_ringoscillator_n5782, inverseur_n227_ringoscillator_n5778, inverseur_n226_ringoscillator_n5774, inverseur_n225_ringoscillator_n5770, inverseur_n224_ringoscillator_n5766, inverseur_n223_ringoscillator_n5762, inverseur_n222_ringoscillator_n5758, inverseur_n221_ringoscillator_n5754, inverseur_n220_ringoscillator_n5750, inverseur_n219_ringoscillator_n5746, inverseur_n218_ringoscillator_n5742, inverseur_n217_ringoscillator_n5738, inverseur_n216_ringoscillator_n5734, inverseur_n215_ringoscillator_n5730, inverseur_n214_ringoscillator_n5726, inverseur_n213_ringoscillator_n5722, inverseur_n212_ringoscillator_n5718, inverseur_n211_ringoscillator_n5714, inverseur_n210_ringoscillator_n5710, inverseur_n209_ringoscillator_n5706, inverseur_n208_ringoscillator_n5702, inverseur_n207_ringoscillator_n5698, inverseur_n206_ringoscillator_n5694, inverseur_n205_ringoscillator_n5690, inverseur_n204_ringoscillator_n5686, inverseur_n203_ringoscillator_n5682, inverseur_n202_ringoscillator_n5678, inverseur_n201_ringoscillator_n5674, inverseur_n200_ringoscillator_n5670, inverseur_n199_ringoscillator_n5666, inverseur_n198_ringoscillator_n5662, inverseur_n197_ringoscillator_n5658, inverseur_n196_ringoscillator_n5654, inverseur_n195_ringoscillator_n5650, inverseur_n194_ringoscillator_n5646, inverseur_n193_ringoscillator_n5642, inverseur_n192_ringoscillator_n5638, inverseur_n191_ringoscillator_n5634, inverseur_n190_ringoscillator_n5630, inverseur_n189_ringoscillator_n5626, inverseur_n188_ringoscillator_n5622, inverseur_n187_ringoscillator_n5618, inverseur_n186_ringoscillator_n5614, inverseur_n185_ringoscillator_n5610, inverseur_n184_ringoscillator_n5606, inverseur_n183_ringoscillator_n5602, inverseur_n182_ringoscillator_n5598, inverseur_n181_ringoscillator_n5594, inverseur_n180_ringoscillator_n5590, inverseur_n179_ringoscillator_n5586, inverseur_n178_ringoscillator_n5582, inverseur_n177_ringoscillator_n5578, inverseur_n176_ringoscillator_n5574, inverseur_n175_ringoscillator_n5570, inverseur_n174_ringoscillator_n5566, inverseur_n173_ringoscillator_n5562, inverseur_n172_ringoscillator_n5558, inverseur_n171_ringoscillator_n5554, inverseur_n170_ringoscillator_n5550, inverseur_n169_ringoscillator_n5546, inverseur_n168_ringoscillator_n5542, inverseur_n167_ringoscillator_n5538, inverseur_n166_ringoscillator_n5534, inverseur_n165_ringoscillator_n5530, inverseur_n164_ringoscillator_n5526, inverseur_n163_ringoscillator_n5522, inverseur_n162_ringoscillator_n5518, inverseur_n161_ringoscillator_n5514, inverseur_n160_ringoscillator_n5510, inverseur_n159_ringoscillator_n5506, inverseur_n158_ringoscillator_n5502, inverseur_n157_ringoscillator_n5498, inverseur_n156_ringoscillator_n5494, inverseur_n155_ringoscillator_n5490, inverseur_n154_ringoscillator_n5486, inverseur_n153_ringoscillator_n5482, inverseur_n152_ringoscillator_n5478, inverseur_n151_ringoscillator_n5474, inverseur_n150_ringoscillator_n5470, inverseur_n149_ringoscillator_n5466, inverseur_n148_ringoscillator_n5462, inverseur_n147_ringoscillator_n5458, inverseur_n146_ringoscillator_n5454, inverseur_n145_ringoscillator_n5450, inverseur_n144_ringoscillator_n5446, inverseur_n143_ringoscillator_n5442, inverseur_n142_ringoscillator_n5438, inverseur_n141_ringoscillator_n5434, inverseur_n140_ringoscillator_n5430, inverseur_n139_ringoscillator_n5426, inverseur_n138_ringoscillator_n5422, inverseur_n137_ringoscillator_n5418, inverseur_n136_ringoscillator_n5414, inverseur_n135_ringoscillator_n5410, inverseur_n134_ringoscillator_n5406, inverseur_n133_ringoscillator_n5402, inverseur_n132_ringoscillator_n5398, inverseur_n131_ringoscillator_n5394, inverseur_n130_ringoscillator_n5390, inverseur_n129_ringoscillator_n5386, inverseur_n128_ringoscillator_n5382, inverseur_n127_ringoscillator_n5378, inverseur_n126_ringoscillator_n5374, inverseur_n125_ringoscillator_n5370, inverseur_n124_ringoscillator_n5366, inverseur_n123_ringoscillator_n5362, inverseur_n122_ringoscillator_n5358, inverseur_n121_ringoscillator_n5354, inverseur_n120_ringoscillator_n5350, inverseur_n119_ringoscillator_n5346, inverseur_n118_ringoscillator_n5342, inverseur_n117_ringoscillator_n5338, inverseur_n116_ringoscillator_n5334, inverseur_n115_ringoscillator_n5330, inverseur_n114_ringoscillator_n5326, inverseur_n113_ringoscillator_n5322, inverseur_n112_ringoscillator_n5318, inverseur_n111_ringoscillator_n5314, inverseur_n110_ringoscillator_n5310, inverseur_n109_ringoscillator_n5306, inverseur_n108_ringoscillator_n5302, inverseur_n107_ringoscillator_n5298, inverseur_n106_ringoscillator_n5294, inverseur_n105_ringoscillator_n5290, inverseur_n104_ringoscillator_n5286, inverseur_n103_ringoscillator_n5282, inverseur_n102_ringoscillator_n5278, inverseur_n101_ringoscillator_n5274, inverseur_n100_ringoscillator_n5270, inverseur_n99_ringoscillator_n5266, inverseur_n98_ringoscillator_n5262, inverseur_n97_ringoscillator_n5258, inverseur_n96_ringoscillator_n5254, inverseur_n95_ringoscillator_n5250, inverseur_n94_ringoscillator_n5246, inverseur_n93_ringoscillator_n5242, inverseur_n92_ringoscillator_n5238, inverseur_n91_ringoscillator_n5234, inverseur_n90_ringoscillator_n5230, inverseur_n89_ringoscillator_n5226, inverseur_n88_ringoscillator_n5222, inverseur_n87_ringoscillator_n5218, inverseur_n86_ringoscillator_n5214, inverseur_n85_ringoscillator_n5210, inverseur_n84_ringoscillator_n5206, inverseur_n83_ringoscillator_n5202, inverseur_n82_ringoscillator_n5198, inverseur_n81_ringoscillator_n5194, inverseur_n80_ringoscillator_n5190, inverseur_n79_ringoscillator_n5186, inverseur_n78_ringoscillator_n5182, inverseur_n77_ringoscillator_n5178, inverseur_n76_ringoscillator_n5174, inverseur_n75_ringoscillator_n5170, inverseur_n74_ringoscillator_n5166, inverseur_n73_ringoscillator_n5162, inverseur_n72_ringoscillator_n5158, inverseur_n71_ringoscillator_n5154, inverseur_n70_ringoscillator_n5150, inverseur_n69_ringoscillator_n5146, inverseur_n68_ringoscillator_n5142, inverseur_n67_ringoscillator_n5138, inverseur_n66_ringoscillator_n5134, inverseur_n65_ringoscillator_n5130, inverseur_n64_ringoscillator_n5126, inverseur_n63_ringoscillator_n5122, inverseur_n62_ringoscillator_n5118, inverseur_n61_ringoscillator_n5114, inverseur_n60_ringoscillator_n5110, inverseur_n59_ringoscillator_n5106, inverseur_n58_ringoscillator_n5102, inverseur_n57_ringoscillator_n5098, inverseur_n56_ringoscillator_n5094, inverseur_n55_ringoscillator_n5090, inverseur_n54_ringoscillator_n5086, inverseur_n53_ringoscillator_n5082, inverseur_n52_ringoscillator_n5078, inverseur_n51_ringoscillator_n5074, inverseur_n50_ringoscillator_n5070, inverseur_n49_ringoscillator_n5066, inverseur_n48_ringoscillator_n5062, inverseur_n47_ringoscillator_n5058, inverseur_n46_ringoscillator_n5054, inverseur_n45_ringoscillator_n5050, inverseur_n44_ringoscillator_n5046, inverseur_n43_ringoscillator_n5042, inverseur_n42_ringoscillator_n5038, inverseur_n41_ringoscillator_n5034, inverseur_n40_ringoscillator_n5030, inverseur_n39_ringoscillator_n5026, inverseur_n38_ringoscillator_n5022, inverseur_n37_ringoscillator_n5018, inverseur_n36_ringoscillator_n5014, inverseur_n35_ringoscillator_n5010, inverseur_n34_ringoscillator_n5006, inverseur_n33_ringoscillator_n5002, inverseur_n32_ringoscillator_n4998, inverseur_n31_ringoscillator_n4994, inverseur_n30_ringoscillator_n4990, inverseur_n29_ringoscillator_n4986, inverseur_n28_ringoscillator_n4982, inverseur_n27_ringoscillator_n4978, inverseur_n26_ringoscillator_n4974, inverseur_n25_ringoscillator_n4970, inverseur_n24_ringoscillator_n4966, inverseur_n23_ringoscillator_n4962, inverseur_n22_ringoscillator_n4958, inverseur_n21_ringoscillator_n4954, inverseur_n20_ringoscillator_n4950, inverseur_n19_ringoscillator_n4946, inverseur_n18_ringoscillator_n4942, inverseur_n17_ringoscillator_n4938, inverseur_n16_ringoscillator_n4934, inverseur_n15_ringoscillator_n4930, inverseur_n14_ringoscillator_n4926, inverseur_n13_ringoscillator_n4922, inverseur_n12_ringoscillator_n4918, inverseur_n11_ringoscillator_n4914, inverseur_n10_ringoscillator_n4910, inverseur_n9_ringoscillator_n4906, inverseur_n8_ringoscillator_n4902, inverseur_n7_ringoscillator_n4898, inverseur_n6_ringoscillator_n4894, inverseur_n5_ringoscillator_n4890, inverseur_n4_ringoscillator_n4886, inverseur_n3_ringoscillator_n4882, inverseur_n2_ringoscillator_n4878, inverseur_n1_ringoscillator_n4874};
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10766_o = n5902_o | n5929_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10767_o = n10766_o | n5947_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10768_o = n10767_o | n5965_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10769_o = n10768_o | n5983_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10770_o = n10769_o | n6001_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10771_o = n10770_o | n6019_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10772_o = n10771_o | n6037_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10773_o = n10772_o | n6055_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10774_o = n10773_o | n6073_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10775_o = n10774_o | n6091_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10776_o = n10775_o | n6109_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10777_o = n10776_o | n6127_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10778_o = n10777_o | n6145_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10779_o = n10778_o | n6163_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10780_o = n10779_o | n6181_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10781_o = n10780_o | n6199_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10782_o = n10781_o | n6217_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10783_o = n10782_o | n6235_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10784_o = n10783_o | n6253_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10785_o = n10784_o | n6271_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10786_o = n10785_o | n6289_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10787_o = n10786_o | n6307_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10788_o = n10787_o | n6325_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10789_o = n10788_o | n6343_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10790_o = n10789_o | n6361_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10791_o = n10790_o | n6379_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10792_o = n10791_o | n6397_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10793_o = n10792_o | n6415_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10794_o = n10793_o | n6433_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10795_o = n10794_o | n6451_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10796_o = n10795_o | n6469_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10797_o = n10796_o | n6487_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10798_o = n10797_o | n6505_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10799_o = n10798_o | n6523_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10800_o = n10799_o | n6541_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10801_o = n10800_o | n6559_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10802_o = n10801_o | n6577_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10803_o = n10802_o | n6595_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10804_o = n10803_o | n6613_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10805_o = n10804_o | n6631_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10806_o = n10805_o | n6649_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10807_o = n10806_o | n6667_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10808_o = n10807_o | n6685_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10809_o = n10808_o | n6703_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10810_o = n10809_o | n6721_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10811_o = n10810_o | n6739_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10812_o = n10811_o | n6757_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10813_o = n10812_o | n6775_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10814_o = n10813_o | n6793_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10815_o = n10814_o | n6811_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10816_o = n10815_o | n6829_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10817_o = n10816_o | n6847_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10818_o = n10817_o | n6865_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10819_o = n10818_o | n6883_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10820_o = n10819_o | n6901_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10821_o = n10820_o | n6919_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10822_o = n10821_o | n6937_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10823_o = n10822_o | n6955_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10824_o = n10823_o | n6973_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10825_o = n10824_o | n6991_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10826_o = n10825_o | n7009_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10827_o = n10826_o | n7027_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10828_o = n10827_o | n7045_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10829_o = n10828_o | n7063_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10830_o = n10829_o | n7081_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10831_o = n10830_o | n7099_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10832_o = n10831_o | n7117_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10833_o = n10832_o | n7135_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10834_o = n10833_o | n7153_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10835_o = n10834_o | n7171_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10836_o = n10835_o | n7189_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10837_o = n10836_o | n7207_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10838_o = n10837_o | n7225_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10839_o = n10838_o | n7243_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10840_o = n10839_o | n7261_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10841_o = n10840_o | n7279_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10842_o = n10841_o | n7297_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10843_o = n10842_o | n7315_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10844_o = n10843_o | n7333_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10845_o = n10844_o | n7351_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10846_o = n10845_o | n7369_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10847_o = n10846_o | n7387_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10848_o = n10847_o | n7405_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10849_o = n10848_o | n7423_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10850_o = n10849_o | n7441_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10851_o = n10850_o | n7459_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10852_o = n10851_o | n7477_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10853_o = n10852_o | n7495_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10854_o = n10853_o | n7513_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10855_o = n10854_o | n7531_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10856_o = n10855_o | n7549_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10857_o = n10856_o | n7567_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10858_o = n10857_o | n7585_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10859_o = n10858_o | n7603_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10860_o = n10859_o | n7621_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10861_o = n10860_o | n7639_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10862_o = n10861_o | n7657_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10863_o = n10862_o | n7675_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10864_o = n10863_o | n7693_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10865_o = n10864_o | n7711_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10866_o = n10865_o | n7729_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10867_o = n10866_o | n7747_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10868_o = n10867_o | n7765_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10869_o = n10868_o | n7783_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10870_o = n10869_o | n7801_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10871_o = n10870_o | n7819_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10872_o = n10871_o | n7837_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10873_o = n10872_o | n7855_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10874_o = n10873_o | n7873_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10875_o = n10874_o | n7891_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10876_o = n10875_o | n7909_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10877_o = n10876_o | n7927_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10878_o = n10877_o | n7945_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10879_o = n10878_o | n7963_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10880_o = n10879_o | n7981_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10881_o = n10880_o | n7999_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10882_o = n10881_o | n8017_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10883_o = n10882_o | n8035_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10884_o = n10883_o | n8053_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10885_o = n10884_o | n8071_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10886_o = n10885_o | n8089_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10887_o = n10886_o | n8107_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10888_o = n10887_o | n8125_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10889_o = n10888_o | n8143_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10890_o = n10889_o | n8161_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10891_o = n10890_o | n8179_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10892_o = n10891_o | n8197_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10893_o = n10892_o | n8215_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10894_o = n10893_o | n8233_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10895_o = n10894_o | n8251_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10896_o = n10895_o | n8269_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10897_o = n10896_o | n8287_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10898_o = n10897_o | n8305_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10899_o = n10898_o | n8323_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10900_o = n10899_o | n8341_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10901_o = n10900_o | n8359_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10902_o = n10901_o | n8377_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10903_o = n10902_o | n8395_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10904_o = n10903_o | n8413_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10905_o = n10904_o | n8431_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10906_o = n10905_o | n8449_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10907_o = n10906_o | n8467_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10908_o = n10907_o | n8485_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10909_o = n10908_o | n8503_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10910_o = n10909_o | n8521_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10911_o = n10910_o | n8539_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10912_o = n10911_o | n8557_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10913_o = n10912_o | n8575_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10914_o = n10913_o | n8593_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10915_o = n10914_o | n8611_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10916_o = n10915_o | n8629_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10917_o = n10916_o | n8647_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10918_o = n10917_o | n8665_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10919_o = n10918_o | n8683_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10920_o = n10919_o | n8701_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10921_o = n10920_o | n8719_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10922_o = n10921_o | n8737_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10923_o = n10922_o | n8755_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10924_o = n10923_o | n8773_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10925_o = n10924_o | n8791_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10926_o = n10925_o | n8809_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10927_o = n10926_o | n8827_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10928_o = n10927_o | n8845_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10929_o = n10928_o | n8863_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10930_o = n10929_o | n8881_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10931_o = n10930_o | n8899_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10932_o = n10931_o | n8917_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10933_o = n10932_o | n8935_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10934_o = n10933_o | n8953_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10935_o = n10934_o | n8971_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10936_o = n10935_o | n8989_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10937_o = n10936_o | n9007_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10938_o = n10937_o | n9025_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10939_o = n10938_o | n9043_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10940_o = n10939_o | n9061_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10941_o = n10940_o | n9079_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10942_o = n10941_o | n9097_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10943_o = n10942_o | n9115_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10944_o = n10943_o | n9133_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10945_o = n10944_o | n9151_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10946_o = n10945_o | n9169_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10947_o = n10946_o | n9187_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10948_o = n10947_o | n9205_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10949_o = n10948_o | n9223_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10950_o = n10949_o | n9241_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10951_o = n10950_o | n9259_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10952_o = n10951_o | n9277_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10953_o = n10952_o | n9295_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10954_o = n10953_o | n9313_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10955_o = n10954_o | n9331_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10956_o = n10955_o | n9349_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10957_o = n10956_o | n9367_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10958_o = n10957_o | n9385_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10959_o = n10958_o | n9403_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10960_o = n10959_o | n9421_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10961_o = n10960_o | n9439_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10962_o = n10961_o | n9457_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10963_o = n10962_o | n9475_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10964_o = n10963_o | n9493_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10965_o = n10964_o | n9511_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10966_o = n10965_o | n9529_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10967_o = n10966_o | n9547_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10968_o = n10967_o | n9565_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10969_o = n10968_o | n9583_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10970_o = n10969_o | n9601_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10971_o = n10970_o | n9619_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10972_o = n10971_o | n9637_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10973_o = n10972_o | n9655_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10974_o = n10973_o | n9673_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10975_o = n10974_o | n9691_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10976_o = n10975_o | n9709_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10977_o = n10976_o | n9727_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10978_o = n10977_o | n9745_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10979_o = n10978_o | n9763_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10980_o = n10979_o | n9781_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10981_o = n10980_o | n9799_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10982_o = n10981_o | n9817_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10983_o = n10982_o | n9835_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10984_o = n10983_o | n9853_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10985_o = n10984_o | n9871_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10986_o = n10985_o | n9889_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10987_o = n10986_o | n9907_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10988_o = n10987_o | n9925_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10989_o = n10988_o | n9943_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10990_o = n10989_o | n9961_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10991_o = n10990_o | n9979_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10992_o = n10991_o | n9997_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10993_o = n10992_o | n10015_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10994_o = n10993_o | n10033_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10995_o = n10994_o | n10051_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10996_o = n10995_o | n10069_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10997_o = n10996_o | n10087_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10998_o = n10997_o | n10105_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n10999_o = n10998_o | n10123_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n11000_o = n10999_o | n10141_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n11001_o = n11000_o | n10159_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n11002_o = n11001_o | n10177_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n11003_o = n11002_o | n10195_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n11004_o = n11003_o | n10213_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n11005_o = n11004_o | n10231_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n11006_o = n11005_o | n10249_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n11007_o = n11006_o | n10267_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n11008_o = n11007_o | n10285_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n11009_o = n11008_o | n10303_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n11010_o = n11009_o | n10321_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n11011_o = n11010_o | n10339_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n11012_o = n11011_o | n10357_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n11013_o = n11012_o | n10375_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n11014_o = n11013_o | n10393_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n11015_o = n11014_o | n10411_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n11016_o = n11015_o | n10429_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n11017_o = n11016_o | n10447_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n11018_o = n11017_o | n10465_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n11019_o = n11018_o | n10483_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n11020_o = n11019_o | n10501_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  assign n11021_o = n11020_o | n10505_o;
  /* RTL_PUF/vhdl/ro_array.vhd:44:1  */
  always @(n11021_o)
    n11022_q <= n10507_o;
endmodule

module uart_tx
  (input  clk,
   input  reset,
   input  [7:0] data_in,
   input  en,
   output busy_out,
   output tx_out);
  (* KEEP="TRUE" *) reg [10:0] cnt;
  (* KEEP="TRUE" *) reg busy;
  (* KEEP="TRUE" *) reg [3:0] bitcnt;
  (* KEEP="TRUE" *) wire n4788_o;
  (* KEEP="TRUE" *) wire n4791_o;
  (* KEEP="TRUE" *) wire [10:0] n4793_o;
  (* KEEP="TRUE" *) wire n4795_o;
  (* KEEP="TRUE" *) wire [3:0] n4797_o;
  (* KEEP="TRUE" *) wire n4801_o;
  (* KEEP="TRUE" *) wire n4803_o;
  (* KEEP="TRUE" *) wire n4805_o;
  (* KEEP="TRUE" *) wire n4806_o;
  (* KEEP="TRUE" *) wire [31:0] n4807_o;
  (* KEEP="TRUE" *) wire [31:0] n4809_o;
  (* KEEP="TRUE" *) wire [2:0] n4810_o;
  (* KEEP="TRUE" *) wire n4814_o;
  (* KEEP="TRUE" *) wire n4816_o;
  (* KEEP="TRUE" *) wire [31:0] n4817_o;
  (* KEEP="TRUE" *) wire n4819_o;
  (* KEEP="TRUE" *) wire n4821_o;
  (* KEEP="TRUE" *) wire [3:0] n4823_o;
  (* KEEP="TRUE" *) wire n4825_o;
  (* KEEP="TRUE" *) wire [10:0] n4828_o;
  (* KEEP="TRUE" *) wire [10:0] n4829_o;
  (* KEEP="TRUE" *) wire n4831_o;
  (* KEEP="TRUE" *) wire [3:0] n4833_o;
  (* KEEP="TRUE" *) wire [31:0] n4834_o;
  (* KEEP="TRUE" *) wire [31:0] n4836_o;
  (* KEEP="TRUE" *) wire [10:0] n4837_o;
  (* KEEP="TRUE" *) wire [10:0] n4838_o;
  (* KEEP="TRUE" *) wire n4839_o;
  (* KEEP="TRUE" *) wire [3:0] n4840_o;
  (* KEEP="TRUE" *) wire n4841_o;
  (* KEEP="TRUE" *) wire [10:0] n4842_o;
  (* KEEP="TRUE" *) wire n4843_o;
  (* KEEP="TRUE" *) wire [3:0] n4844_o;
  (* KEEP="TRUE" *) reg [10:0] n4852_q;
  (* KEEP="TRUE" *) reg n4853_q;
  (* KEEP="TRUE" *) reg [3:0] n4854_q;
  (* KEEP="TRUE" *) reg n4857_q;
  (* KEEP="TRUE" *) wire n4858_o;
  (* KEEP="TRUE" *) wire n4859_o;
  (* KEEP="TRUE" *) wire n4860_o;
  (* KEEP="TRUE" *) wire n4861_o;
  (* KEEP="TRUE" *) wire n4862_o;
  (* KEEP="TRUE" *) wire n4863_o;
  (* KEEP="TRUE" *) wire n4864_o;
  (* KEEP="TRUE" *) wire n4865_o;
  (* KEEP="TRUE" *) wire [1:0] n4866_o;
  (* KEEP="TRUE" *) reg n4867_o;
  (* KEEP="TRUE" *) wire [1:0] n4868_o;
  (* KEEP="TRUE" *) reg n4869_o;
  (* KEEP="TRUE" *) wire n4870_o;
  (* KEEP="TRUE" *) wire n4871_o;
  assign busy_out = busy;
  assign tx_out = n4857_q;
  /* RTL_PUF/vhdl/UART_TX.vhd:19:12  */
  always @*
    cnt = n4852_q; // (isignal)
  initial
    cnt = 11'b00000000000;
  /* RTL_PUF/vhdl/UART_TX.vhd:20:12  */
  always @*
    busy = n4853_q; // (isignal)
  initial
    busy = 1'b1;
  /* RTL_PUF/vhdl/UART_TX.vhd:21:12  */
  always @*
    bitcnt = n4854_q; // (isignal)
  initial
    bitcnt = 4'b0000;
  /* RTL_PUF/vhdl/UART_TX.vhd:32:13  */
  assign n4788_o = ~busy;
  /* RTL_PUF/vhdl/UART_TX.vhd:33:9  */
  assign n4791_o = en ? 1'b0 : 1'b1;
  /* RTL_PUF/vhdl/UART_TX.vhd:33:9  */
  assign n4793_o = en ? 11'b10011100001 : cnt;
  /* RTL_PUF/vhdl/UART_TX.vhd:33:9  */
  assign n4795_o = en ? 1'b1 : busy;
  /* RTL_PUF/vhdl/UART_TX.vhd:33:9  */
  assign n4797_o = en ? 4'b0000 : bitcnt;
  /* RTL_PUF/vhdl/UART_TX.vhd:46:19  */
  assign n4801_o = bitcnt == 4'b0000;
  /* RTL_PUF/vhdl/UART_TX.vhd:48:22  */
  assign n4803_o = $unsigned(bitcnt) >= $unsigned(4'b0001);
  /* RTL_PUF/vhdl/UART_TX.vhd:48:38  */
  assign n4805_o = $unsigned(bitcnt) < $unsigned(4'b1001);
  /* RTL_PUF/vhdl/UART_TX.vhd:48:27  */
  assign n4806_o = n4805_o & n4803_o;
  /* RTL_PUF/vhdl/UART_TX.vhd:49:31  */
  assign n4807_o = {28'b0, bitcnt};  //  uext
  /* RTL_PUF/vhdl/UART_TX.vhd:49:51  */
  assign n4809_o = n4807_o - 32'b00000000000000000000000000000001;
  /* RTL_PUF/vhdl/UART_TX.vhd:49:51  */
  assign n4810_o = n4809_o[2:0];  // trunc
  /* RTL_PUF/vhdl/UART_TX.vhd:48:9  */
  assign n4814_o = n4806_o ? n4871_o : 1'b1;
  /* RTL_PUF/vhdl/UART_TX.vhd:46:9  */
  assign n4816_o = n4801_o ? 1'b0 : n4814_o;
  /* RTL_PUF/vhdl/UART_TX.vhd:54:16  */
  assign n4817_o = {21'b0, cnt};  //  uext
  /* RTL_PUF/vhdl/UART_TX.vhd:54:16  */
  assign n4819_o = n4817_o == 32'b00000000000000000000000000000000;
  /* RTL_PUF/vhdl/UART_TX.vhd:55:23  */
  assign n4821_o = $unsigned(bitcnt) < $unsigned(4'b1001);
  /* RTL_PUF/vhdl/UART_TX.vhd:56:34  */
  assign n4823_o = bitcnt + 4'b0001;
  /* RTL_PUF/vhdl/UART_TX.vhd:57:27  */
  assign n4825_o = $unsigned(bitcnt) < $unsigned(4'b1000);
  /* RTL_PUF/vhdl/UART_TX.vhd:57:17  */
  assign n4828_o = n4825_o ? 11'b10011100001 : 11'b10001111110;
  /* RTL_PUF/vhdl/UART_TX.vhd:55:13  */
  assign n4829_o = n4821_o ? n4828_o : cnt;
  /* RTL_PUF/vhdl/UART_TX.vhd:55:13  */
  assign n4831_o = n4821_o ? busy : 1'b0;
  /* RTL_PUF/vhdl/UART_TX.vhd:55:13  */
  assign n4833_o = n4821_o ? n4823_o : 4'b0000;
  /* RTL_PUF/vhdl/UART_TX.vhd:68:24  */
  assign n4834_o = {21'b0, cnt};  //  uext
  /* RTL_PUF/vhdl/UART_TX.vhd:68:24  */
  assign n4836_o = n4834_o - 32'b00000000000000000000000000000001;
  /* RTL_PUF/vhdl/UART_TX.vhd:68:20  */
  assign n4837_o = n4836_o[10:0];  // trunc
  /* RTL_PUF/vhdl/UART_TX.vhd:54:9  */
  assign n4838_o = n4819_o ? n4829_o : n4837_o;
  /* RTL_PUF/vhdl/UART_TX.vhd:54:9  */
  assign n4839_o = n4819_o ? n4831_o : busy;
  /* RTL_PUF/vhdl/UART_TX.vhd:54:9  */
  assign n4840_o = n4819_o ? n4833_o : bitcnt;
  /* RTL_PUF/vhdl/UART_TX.vhd:32:5  */
  assign n4841_o = n4788_o ? n4791_o : n4816_o;
  /* RTL_PUF/vhdl/UART_TX.vhd:32:5  */
  assign n4842_o = n4788_o ? n4793_o : n4838_o;
  /* RTL_PUF/vhdl/UART_TX.vhd:32:5  */
  assign n4843_o = n4788_o ? n4795_o : n4839_o;
  /* RTL_PUF/vhdl/UART_TX.vhd:32:5  */
  assign n4844_o = n4788_o ? n4797_o : n4840_o;
  /* RTL_PUF/vhdl/UART_TX.vhd:29:1  */
  always @(posedge clk)
    n4852_q <= n4842_o;
  initial
    n4852_q = 11'b00000000000;
  /* RTL_PUF/vhdl/UART_TX.vhd:29:1  */
  always @(posedge clk)
    n4853_q <= n4843_o;
  initial
    n4853_q = 1'b1;
  /* RTL_PUF/vhdl/UART_TX.vhd:29:1  */
  always @(posedge clk)
    n4854_q <= n4844_o;
  initial
    n4854_q = 4'b0000;
  /* RTL_PUF/vhdl/UART_TX.vhd:29:1  */
  always @(posedge clk)
    n4857_q <= n4841_o;
  /* RTL_PUF/vhdl/UART_TX.vhd:11:8  */
  assign n4858_o = data_in[0];
  /* RTL_PUF/vhdl/UART_TX.vhd:10:8  */
  assign n4859_o = data_in[1];
  /* RTL_PUF/vhdl/UART_TX.vhd:29:1  */
  assign n4860_o = data_in[2];
  /* RTL_PUF/vhdl/UART_TX.vhd:29:1  */
  assign n4861_o = data_in[3];
  assign n4862_o = data_in[4];
  /* RTL_PUF/vhdl/UART_TX.vhd:29:1  */
  assign n4863_o = data_in[5];
  /* RTL_PUF/vhdl/UART_TX.vhd:32:5  */
  assign n4864_o = data_in[6];
  assign n4865_o = data_in[7];
  /* RTL_PUF/vhdl/UART_TX.vhd:49:30  */
  assign n4866_o = n4810_o[1:0];
  /* RTL_PUF/vhdl/UART_TX.vhd:49:30  */
  always @*
    case (n4866_o)
      2'b00: n4867_o = n4858_o;
      2'b01: n4867_o = n4859_o;
      2'b10: n4867_o = n4860_o;
      2'b11: n4867_o = n4861_o;
    endcase
  /* RTL_PUF/vhdl/UART_TX.vhd:49:30  */
  assign n4868_o = n4810_o[1:0];
  /* RTL_PUF/vhdl/UART_TX.vhd:49:30  */
  always @*
    case (n4868_o)
      2'b00: n4869_o = n4862_o;
      2'b01: n4869_o = n4863_o;
      2'b10: n4869_o = n4864_o;
      2'b11: n4869_o = n4865_o;
    endcase
  /* RTL_PUF/vhdl/UART_TX.vhd:49:30  */
  assign n4870_o = n4810_o[2];
  /* RTL_PUF/vhdl/UART_TX.vhd:49:30  */
  assign n4871_o = n4870_o ? n4869_o : n4867_o;
endmodule

module uart_rx
  (input  clk,
   input  rx_in,
   output busy_out,
   output rdy,
   output [7:0] data_out);
  (* KEEP="TRUE" *) reg [10:0] cnt;
  (* KEEP="TRUE" *) reg rx_data;
  (* KEEP="TRUE" *) reg busy;
  (* KEEP="TRUE" *) reg [3:0] num_bits;
  (* KEEP="TRUE" *) reg [7:0] data_out_buf;
  (* KEEP="TRUE" *) wire n4656_o;
  (* KEEP="TRUE" *) wire n4657_o;
  (* KEEP="TRUE" *) wire n4659_o;
  (* KEEP="TRUE" *) wire [3:0] n4661_o;
  (* KEEP="TRUE" *) wire [31:0] n4662_o;
  (* KEEP="TRUE" *) wire n4664_o;
  (* KEEP="TRUE" *) wire n4666_o;
  (* KEEP="TRUE" *) wire n4667_o;
  (* KEEP="TRUE" *) wire [3:0] n4669_o;
  (* KEEP="TRUE" *) wire n4671_o;
  (* KEEP="TRUE" *) wire [31:0] n4672_o;
  (* KEEP="TRUE" *) wire [31:0] n4674_o;
  (* KEEP="TRUE" *) wire [2:0] n4675_o;
  (* KEEP="TRUE" *) wire [3:0] n4679_o;
  (* KEEP="TRUE" *) wire n4681_o;
  (* KEEP="TRUE" *) wire [7:0] n4682_o;
  (* KEEP="TRUE" *) wire n4685_o;
  (* KEEP="TRUE" *) wire [3:0] n4686_o;
  (* KEEP="TRUE" *) wire n4688_o;
  (* KEEP="TRUE" *) wire [7:0] n4689_o;
  (* KEEP="TRUE" *) wire n4690_o;
  (* KEEP="TRUE" *) wire [3:0] n4691_o;
  (* KEEP="TRUE" *) wire [31:0] n4693_o;
  (* KEEP="TRUE" *) wire [31:0] n4695_o;
  (* KEEP="TRUE" *) wire [10:0] n4696_o;
  (* KEEP="TRUE" *) wire n4697_o;
  (* KEEP="TRUE" *) wire [7:0] n4698_o;
  (* KEEP="TRUE" *) wire [10:0] n4700_o;
  (* KEEP="TRUE" *) wire n4701_o;
  (* KEEP="TRUE" *) wire [3:0] n4702_o;
  (* KEEP="TRUE" *) wire n4705_o;
  (* KEEP="TRUE" *) wire [7:0] n4706_o;
  (* KEEP="TRUE" *) wire [10:0] n4708_o;
  (* KEEP="TRUE" *) wire n4709_o;
  (* KEEP="TRUE" *) wire [3:0] n4710_o;
  (* KEEP="TRUE" *) reg [10:0] n4721_q;
  (* KEEP="TRUE" *) reg n4722_q;
  (* KEEP="TRUE" *) reg n4723_q;
  (* KEEP="TRUE" *) reg [3:0] n4724_q;
  (* KEEP="TRUE" *) wire n4725_o;
  (* KEEP="TRUE" *) wire n4726_o;
  (* KEEP="TRUE" *) wire n4727_o;
  (* KEEP="TRUE" *) wire n4728_o;
  (* KEEP="TRUE" *) wire n4729_o;
  (* KEEP="TRUE" *) wire n4730_o;
  (* KEEP="TRUE" *) reg [7:0] n4732_q;
  (* KEEP="TRUE" *) reg n4733_q;
  (* KEEP="TRUE" *) reg n4734_q;
  (* KEEP="TRUE" *) reg [7:0] n4735_q;
  (* KEEP="TRUE" *) wire n4736_o;
  (* KEEP="TRUE" *) wire n4737_o;
  (* KEEP="TRUE" *) wire n4738_o;
  (* KEEP="TRUE" *) wire n4739_o;
  (* KEEP="TRUE" *) wire n4740_o;
  (* KEEP="TRUE" *) wire n4741_o;
  (* KEEP="TRUE" *) wire n4742_o;
  (* KEEP="TRUE" *) wire n4743_o;
  (* KEEP="TRUE" *) wire n4744_o;
  (* KEEP="TRUE" *) wire n4745_o;
  (* KEEP="TRUE" *) wire n4746_o;
  (* KEEP="TRUE" *) wire n4747_o;
  (* KEEP="TRUE" *) wire n4748_o;
  (* KEEP="TRUE" *) wire n4749_o;
  (* KEEP="TRUE" *) wire n4750_o;
  (* KEEP="TRUE" *) wire n4751_o;
  (* KEEP="TRUE" *) wire n4752_o;
  (* KEEP="TRUE" *) wire n4753_o;
  (* KEEP="TRUE" *) wire n4754_o;
  (* KEEP="TRUE" *) wire n4755_o;
  (* KEEP="TRUE" *) wire n4756_o;
  (* KEEP="TRUE" *) wire n4757_o;
  (* KEEP="TRUE" *) wire n4758_o;
  (* KEEP="TRUE" *) wire n4759_o;
  (* KEEP="TRUE" *) wire n4760_o;
  (* KEEP="TRUE" *) wire n4761_o;
  (* KEEP="TRUE" *) wire n4762_o;
  (* KEEP="TRUE" *) wire n4763_o;
  (* KEEP="TRUE" *) wire n4764_o;
  (* KEEP="TRUE" *) wire n4765_o;
  (* KEEP="TRUE" *) wire n4766_o;
  (* KEEP="TRUE" *) wire n4767_o;
  (* KEEP="TRUE" *) wire n4768_o;
  (* KEEP="TRUE" *) wire n4769_o;
  (* KEEP="TRUE" *) wire n4770_o;
  (* KEEP="TRUE" *) wire n4771_o;
  (* KEEP="TRUE" *) wire n4772_o;
  (* KEEP="TRUE" *) wire n4773_o;
  (* KEEP="TRUE" *) wire n4774_o;
  (* KEEP="TRUE" *) wire n4775_o;
  (* KEEP="TRUE" *) wire n4776_o;
  (* KEEP="TRUE" *) wire n4777_o;
  (* KEEP="TRUE" *) wire [7:0] n4778_o;
  assign busy_out = n4733_q;
  assign rdy = n4734_q;
  assign data_out = n4735_q;
  /* RTL_PUF/vhdl/UART_RX.vhd:18:12  */
  always @*
    cnt = n4721_q; // (isignal)
  initial
    cnt = 11'b00000000000;
  /* RTL_PUF/vhdl/UART_RX.vhd:19:12  */
  always @*
    rx_data = n4722_q; // (isignal)
  initial
    rx_data = 1'b0;
  /* RTL_PUF/vhdl/UART_RX.vhd:20:12  */
  always @*
    busy = n4723_q; // (isignal)
  initial
    busy = 1'b0;
  /* RTL_PUF/vhdl/UART_RX.vhd:21:12  */
  always @*
    num_bits = n4724_q; // (isignal)
  initial
    num_bits = 4'b0000;
  /* RTL_PUF/vhdl/UART_RX.vhd:22:12  */
  always @*
    data_out_buf = n4732_q; // (isignal)
  initial
    data_out_buf = 8'b00000000;
  /* RTL_PUF/vhdl/UART_RX.vhd:35:13  */
  assign n4656_o = ~busy;
  /* RTL_PUF/vhdl/UART_RX.vhd:37:20  */
  assign n4657_o = ~rx_data;
  /* RTL_PUF/vhdl/UART_RX.vhd:37:9  */
  assign n4659_o = n4657_o ? 1'b1 : busy;
  /* RTL_PUF/vhdl/UART_RX.vhd:37:9  */
  assign n4661_o = n4657_o ? 4'b0000 : num_bits;
  /* RTL_PUF/vhdl/UART_RX.vhd:48:16  */
  assign n4662_o = {21'b0, cnt};  //  uext
  /* RTL_PUF/vhdl/UART_RX.vhd:48:16  */
  assign n4664_o = n4662_o == 32'b00000000000000000000000000000000;
  /* RTL_PUF/vhdl/UART_RX.vhd:50:25  */
  assign n4666_o = num_bits == 4'b0000;
  /* RTL_PUF/vhdl/UART_RX.vhd:51:25  */
  assign n4667_o = ~rx_data;
  /* RTL_PUF/vhdl/UART_RX.vhd:52:38  */
  assign n4669_o = num_bits + 4'b0001;
  /* RTL_PUF/vhdl/UART_RX.vhd:53:28  */
  assign n4671_o = num_bits == 4'b1001;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:30  */
  assign n4672_o = {28'b0, num_bits};  //  uext
  /* RTL_PUF/vhdl/UART_RX.vhd:58:52  */
  assign n4674_o = n4672_o - 32'b00000000000000000000000000000001;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:52  */
  assign n4675_o = n4674_o[2:0];  // trunc
  /* RTL_PUF/vhdl/UART_RX.vhd:60:38  */
  assign n4679_o = num_bits + 4'b0001;
  /* RTL_PUF/vhdl/UART_RX.vhd:53:13  */
  assign n4681_o = n4671_o ? 1'b1 : n4734_q;
  /* RTL_PUF/vhdl/UART_RX.vhd:53:13  */
  assign n4682_o = n4671_o ? data_out_buf : n4735_q;
  /* RTL_PUF/vhdl/UART_RX.vhd:53:13  */
  assign n4685_o = n4671_o ? 1'b0 : 1'b1;
  /* RTL_PUF/vhdl/UART_RX.vhd:53:13  */
  assign n4686_o = n4671_o ? num_bits : n4679_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:50:13  */
  assign n4688_o = n4666_o ? n4734_q : n4681_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:50:13  */
  assign n4689_o = n4666_o ? n4735_q : n4682_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:50:13  */
  assign n4690_o = n4666_o ? n4667_o : n4685_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:50:13  */
  assign n4691_o = n4666_o ? n4669_o : n4686_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:66:24  */
  assign n4693_o = {21'b0, cnt};  //  uext
  /* RTL_PUF/vhdl/UART_RX.vhd:66:24  */
  assign n4695_o = n4693_o - 32'b00000000000000000000000000000001;
  /* RTL_PUF/vhdl/UART_RX.vhd:66:20  */
  assign n4696_o = n4695_o[10:0];  // trunc
  /* RTL_PUF/vhdl/UART_RX.vhd:48:9  */
  assign n4697_o = n4664_o ? n4688_o : n4734_q;
  /* RTL_PUF/vhdl/UART_RX.vhd:48:9  */
  assign n4698_o = n4664_o ? n4689_o : n4735_q;
  /* RTL_PUF/vhdl/UART_RX.vhd:48:9  */
  assign n4700_o = n4664_o ? 11'b10011100001 : n4696_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:48:9  */
  assign n4701_o = n4664_o ? n4690_o : busy;
  /* RTL_PUF/vhdl/UART_RX.vhd:48:9  */
  assign n4702_o = n4664_o ? n4691_o : num_bits;
  /* RTL_PUF/vhdl/UART_RX.vhd:35:5  */
  assign n4705_o = n4656_o ? 1'b0 : n4697_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:35:5  */
  assign n4706_o = n4656_o ? n4735_q : n4698_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:35:5  */
  assign n4708_o = n4656_o ? 11'b01001110000 : n4700_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:35:5  */
  assign n4709_o = n4656_o ? n4659_o : n4701_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:35:5  */
  assign n4710_o = n4656_o ? n4661_o : n4702_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:33:1  */
  always @(posedge clk)
    n4721_q <= n4708_o;
  initial
    n4721_q = 11'b00000000000;
  /* RTL_PUF/vhdl/UART_RX.vhd:33:1  */
  always @(posedge clk)
    n4722_q <= rx_in;
  initial
    n4722_q = 1'b0;
  /* RTL_PUF/vhdl/UART_RX.vhd:33:1  */
  always @(posedge clk)
    n4723_q <= n4709_o;
  initial
    n4723_q = 1'b0;
  /* RTL_PUF/vhdl/UART_RX.vhd:33:1  */
  always @(posedge clk)
    n4724_q <= n4710_o;
  initial
    n4724_q = 4'b0000;
  /* RTL_PUF/vhdl/UART_RX.vhd:35:5  */
  assign n4725_o = ~n4656_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:35:5  */
  assign n4726_o = n4725_o & n4664_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:50:13  */
  assign n4727_o = ~n4666_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:35:5  */
  assign n4728_o = n4726_o & n4727_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:53:13  */
  assign n4729_o = ~n4671_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:35:5  */
  assign n4730_o = n4728_o & n4729_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:33:1  */
  always @(posedge clk)
    n4732_q <= n4778_o;
  initial
    n4732_q = 8'b00000000;
  /* RTL_PUF/vhdl/UART_RX.vhd:33:1  */
  always @(posedge clk)
    n4733_q <= busy;
  /* RTL_PUF/vhdl/UART_RX.vhd:33:1  */
  always @(posedge clk)
    n4734_q <= n4705_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:33:1  */
  always @(posedge clk)
    n4735_q <= n4706_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4736_o = n4675_o[2];
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4737_o = ~n4736_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4738_o = n4675_o[1];
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4739_o = ~n4738_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4740_o = n4737_o & n4739_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4741_o = n4737_o & n4738_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4742_o = n4736_o & n4739_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4743_o = n4736_o & n4738_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4744_o = n4675_o[0];
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4745_o = ~n4744_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4746_o = n4740_o & n4745_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4747_o = n4740_o & n4744_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4748_o = n4741_o & n4745_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4749_o = n4741_o & n4744_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4750_o = n4742_o & n4745_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4751_o = n4742_o & n4744_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4752_o = n4743_o & n4745_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4753_o = n4743_o & n4744_o;
  assign n4754_o = data_out_buf[0];
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4755_o = n4746_o & n4730_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4756_o = n4755_o ? rx_data : n4754_o;
  assign n4757_o = data_out_buf[1];
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4758_o = n4747_o & n4730_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4759_o = n4758_o ? rx_data : n4757_o;
  assign n4760_o = data_out_buf[2];
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4761_o = n4748_o & n4730_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4762_o = n4761_o ? rx_data : n4760_o;
  assign n4763_o = data_out_buf[3];
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4764_o = n4749_o & n4730_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4765_o = n4764_o ? rx_data : n4763_o;
  assign n4766_o = data_out_buf[4];
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4767_o = n4750_o & n4730_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4768_o = n4767_o ? rx_data : n4766_o;
  assign n4769_o = data_out_buf[5];
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4770_o = n4751_o & n4730_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4771_o = n4770_o ? rx_data : n4769_o;
  assign n4772_o = data_out_buf[6];
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4773_o = n4752_o & n4730_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4774_o = n4773_o ? rx_data : n4772_o;
  assign n4775_o = data_out_buf[7];
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4776_o = n4753_o & n4730_o;
  /* RTL_PUF/vhdl/UART_RX.vhd:58:17  */
  assign n4777_o = n4776_o ? rx_data : n4775_o;
  assign n4778_o = {n4777_o, n4774_o, n4771_o, n4768_o, n4765_o, n4762_o, n4759_o, n4756_o};
endmodule

module ro_puf_s7
  (input  clk,
   input  uart_rx,
   input  reset_btn,
   output led1,
   output led2,
   output led3,
   output led4,
   output uart_tx,
   output ledR_1,
   output ledG_1,
   output ledB_1);
  (* KEEP="TRUE" *) wire [7:0] received_word;
  (* KEEP="TRUE" *) wire rdy;
  (* KEEP="TRUE" *) reg tx_en;
  (* KEEP="TRUE" *) wire tx_busy;
  (* KEEP="TRUE" *) reg [7:0] tx_data_in;
  (* KEEP="TRUE" *) reg shift_state;
  (* KEEP="TRUE" *) reg [7:0] output_data;
  (* KEEP="TRUE" *) reg [7:0] internal_challenge_mux;
  (* KEEP="TRUE" *) localparam [63:0] n18_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  (* KEEP="TRUE" *) reg [63:0] puf_response;
  (* KEEP="TRUE" *) reg puf_start;
  (* KEEP="TRUE" *) reg [7:0] mux_1_challenge;
  (* KEEP="TRUE" *) reg [7:0] mux_2_challenge;
  (* KEEP="TRUE" *) reg mux_1_out;
  (* KEEP="TRUE" *) reg mux_2_out;
  (* KEEP="TRUE" *) reg [28:0] compteur_cycles;
  (* KEEP="TRUE" *) reg [30:0] mux_1_counter;
  (* KEEP="TRUE" *) reg [30:0] mux_2_counter;
  (* KEEP="TRUE" *) reg [255:0] enable_1;
  (* KEEP="TRUE" *) reg [255:0] enable_2;
  (* KEEP="TRUE" *) reg reset_counter;
  (* KEEP="TRUE" *) reg enable_comparison;
  (* KEEP="TRUE" *) reg enable_counter;
  (* KEEP="TRUE" *) reg data_valid;
  (* KEEP="TRUE" *) reg tx_available;
  (* KEEP="TRUE" *) wire [2:0] counter_timer;
  (* KEEP="TRUE" *) reg [31:0] timer_size;
  (* KEEP="TRUE" *) reg [255:0] ro_filter;
  (* KEEP="TRUE" *) reg [7:0] rom_address;
  (* KEEP="TRUE" *) wire [15:0] rom_data_out;
  (* KEEP="TRUE" *) reg mode_select;
  (* KEEP="TRUE" *) wire [2:0] state;
  (* KEEP="TRUE" *) reg [4:0] transmission_state;
  (* KEEP="TRUE" *) wire uart_rx_inst_busy_out;
  (* KEEP="TRUE" *) wire uart_rx_inst_rdy;
  (* KEEP="TRUE" *) wire [7:0] uart_rx_inst_data_out;
  (* KEEP="TRUE" *) wire uart_tx_inst_busy_out;
  (* KEEP="TRUE" *) wire uart_tx_inst_tx_out;
  (* KEEP="TRUE" *) wire n47_o;
  (* KEEP="TRUE" *) wire [4:0] n50_o;
  (* KEEP="TRUE" *) wire n52_o;
  (* KEEP="TRUE" *) wire [7:0] n53_o;
  (* KEEP="TRUE" *) wire n55_o;
  (* KEEP="TRUE" *) wire n57_o;
  (* KEEP="TRUE" *) wire [7:0] n58_o;
  (* KEEP="TRUE" *) wire n60_o;
  (* KEEP="TRUE" *) wire n62_o;
  (* KEEP="TRUE" *) wire [7:0] n63_o;
  (* KEEP="TRUE" *) wire n65_o;
  (* KEEP="TRUE" *) wire n67_o;
  (* KEEP="TRUE" *) wire [7:0] n68_o;
  (* KEEP="TRUE" *) wire n70_o;
  (* KEEP="TRUE" *) wire n72_o;
  (* KEEP="TRUE" *) wire [7:0] n73_o;
  (* KEEP="TRUE" *) wire n75_o;
  (* KEEP="TRUE" *) wire n77_o;
  (* KEEP="TRUE" *) wire [7:0] n78_o;
  (* KEEP="TRUE" *) wire n80_o;
  (* KEEP="TRUE" *) wire n82_o;
  (* KEEP="TRUE" *) wire [7:0] n83_o;
  (* KEEP="TRUE" *) wire n85_o;
  (* KEEP="TRUE" *) wire n87_o;
  (* KEEP="TRUE" *) wire [7:0] n88_o;
  (* KEEP="TRUE" *) wire n90_o;
  (* KEEP="TRUE" *) wire n92_o;
  (* KEEP="TRUE" *) wire [16:0] n93_o;
  (* KEEP="TRUE" *) reg n111_o;
  (* KEEP="TRUE" *) reg [7:0] n112_o;
  (* KEEP="TRUE" *) reg n115_o;
  (* KEEP="TRUE" *) reg [4:0] n133_o;
  (* KEEP="TRUE" *) wire n146_o;
  (* KEEP="TRUE" *) wire n149_o;
  (* KEEP="TRUE" *) wire n152_o;
  (* KEEP="TRUE" *) wire n154_o;
  (* KEEP="TRUE" *) wire [1:0] n155_o;
  (* KEEP="TRUE" *) reg n159_o;
  (* KEEP="TRUE" *) reg n162_o;
  (* KEEP="TRUE" *) wire [6:0] n163_o;
  (* KEEP="TRUE" *) wire [6:0] n164_o;
  (* KEEP="TRUE" *) reg [6:0] n166_o;
  (* KEEP="TRUE" *) wire n167_o;
  (* KEEP="TRUE" *) reg n169_o;
  (* KEEP="TRUE" *) wire n171_o;
  (* KEEP="TRUE" *) wire n174_o;
  (* KEEP="TRUE" *) wire n176_o;
  (* KEEP="TRUE" *) wire [7:0] n177_o;
  (* KEEP="TRUE" *) wire [7:0] n178_o;
  (* KEEP="TRUE" *) wire n184_o;
  (* KEEP="TRUE" *) wire n185_o;
  (* KEEP="TRUE" *) wire [2:0] n186_o;
  (* KEEP="TRUE" *) localparam n187_o = 1'b0;
  (* KEEP="TRUE" *) localparam n188_o = 1'b0;
  (* KEEP="TRUE" *) wire uut1_n189;
  (* KEEP="TRUE" *) wire uut1_output ;
  (* KEEP="TRUE" *) wire uut2_n192;
  (* KEEP="TRUE" *) wire uut2_output ;
  (* KEEP="TRUE" *) wire [15:0] rom_n195;
  (* KEEP="TRUE" *) wire n201_o;
  (* KEEP="TRUE" *) wire n203_o;
  (* KEEP="TRUE" *) wire n205_o;
  (* KEEP="TRUE" *) wire n207_o;
  (* KEEP="TRUE" *) wire [31:0] n210_o;
  (* KEEP="TRUE" *) wire [31:0] n212_o;
  (* KEEP="TRUE" *) wire [31:0] n214_o;
  (* KEEP="TRUE" *) wire [31:0] n216_o;
  (* KEEP="TRUE" *) wire [28:0] n223_o;
  (* KEEP="TRUE" *) wire [28:0] n225_o;
  (* KEEP="TRUE" *) wire n231_o;
  (* KEEP="TRUE" *) wire [7:0] n232_o;
  (* KEEP="TRUE" *) wire [7:0] n233_o;
  (* KEEP="TRUE" *) wire [7:0] n234_o;
  (* KEEP="TRUE" *) wire [7:0] n235_o;
  (* KEEP="TRUE" *) wire n236_o;
  (* KEEP="TRUE" *) wire [2:0] n242_o;
  (* KEEP="TRUE" *) wire [2:0] n247_o;
  (* KEEP="TRUE" *) wire [2:0] n248_o;
  (* KEEP="TRUE" *) wire [2:0] n250_o;
  (* KEEP="TRUE" *) wire n252_o;
  (* KEEP="TRUE" *) wire n253_o;
  (* KEEP="TRUE" *) wire [7:0] n262_o;
  (* KEEP="TRUE" *) wire [7:0] n267_o;
  (* KEEP="TRUE" *) wire [255:0] n272_o;
  (* KEEP="TRUE" *) wire [255:0] n273_o;
  (* KEEP="TRUE" *) wire [30:0] n274_o;
  (* KEEP="TRUE" *) wire [28:0] n275_o;
  (* KEEP="TRUE" *) wire n276_o;
  (* KEEP="TRUE" *) wire [2:0] n279_o;
  (* KEEP="TRUE" *) wire n281_o;
  (* KEEP="TRUE" *) wire [2:0] n284_o;
  (* KEEP="TRUE" *) wire n286_o;
  (* KEEP="TRUE" *) wire n287_o;
  (* KEEP="TRUE" *) wire n289_o;
  (* KEEP="TRUE" *) wire [2:0] n292_o;
  (* KEEP="TRUE" *) wire [31:0] n293_o;
  (* KEEP="TRUE" *) wire n295_o;
  (* KEEP="TRUE" *) wire [2:0] n298_o;
  (* KEEP="TRUE" *) wire [2:0] n299_o;
  (* KEEP="TRUE" *) wire n301_o;
  (* KEEP="TRUE" *) wire n302_o;
  (* KEEP="TRUE" *) wire [7:0] n304_o;
  (* KEEP="TRUE" *) wire [31:0] n305_o;
  (* KEEP="TRUE" *) wire [31:0] n307_o;
  (* KEEP="TRUE" *) wire [7:0] n308_o;
  (* KEEP="TRUE" *) wire [7:0] n309_o;
  (* KEEP="TRUE" *) wire [7:0] n310_o;
  (* KEEP="TRUE" *) wire n312_o;
  (* KEEP="TRUE" *) wire n313_o;
  (* KEEP="TRUE" *) wire n318_o;
  (* KEEP="TRUE" *) wire [2:0] n321_o;
  (* KEEP="TRUE" *) wire [2:0] n323_o;
  (* KEEP="TRUE" *) wire [31:0] n326_o;
  (* KEEP="TRUE" *) wire n328_o;
  (* KEEP="TRUE" *) wire [2:0] n331_o;
  (* KEEP="TRUE" *) wire [2:0] n333_o;
  (* KEEP="TRUE" *) wire [2:0] n334_o;
  (* KEEP="TRUE" *) wire n336_o;
  (* KEEP="TRUE" *) wire [5:0] n337_o;
  (* KEEP="TRUE" *) reg n344_o;
  (* KEEP="TRUE" *) reg n351_o;
  (* KEEP="TRUE" *) reg n358_o;
  (* KEEP="TRUE" *) reg [7:0] n361_o;
  (* KEEP="TRUE" *) reg [255:0] n365_o;
  (* KEEP="TRUE" *) reg [255:0] n369_o;
  (* KEEP="TRUE" *) reg n376_o;
  (* KEEP="TRUE" *) reg n383_o;
  (* KEEP="TRUE" *) reg n390_o;
  (* KEEP="TRUE" *) reg [7:0] n393_o;
  (* KEEP="TRUE" *) reg [2:0] n396_o;
  (* KEEP="TRUE" *) wire [30:0] n415_o;
  (* KEEP="TRUE" *) wire [30:0] n422_o;
  (* KEEP="TRUE" *) wire n431_o;
  (* KEEP="TRUE" *) wire [61:0] n434_o;
  (* KEEP="TRUE" *) wire [61:0] n435_o;
  (* KEEP="TRUE" *) wire [61:0] n436_o;
  (* KEEP="TRUE" *) wire n437_o;
  (* KEEP="TRUE" *) wire n444_o;
  (* KEEP="TRUE" *) wire n451_o;
  (* KEEP="TRUE" *) reg n452_q;
  (* KEEP="TRUE" *) wire [7:0] n453_o;
  (* KEEP="TRUE" *) reg [7:0] n454_q;
  (* KEEP="TRUE" *) reg n455_q;
  (* KEEP="TRUE" *) reg [7:0] n456_q;
  (* KEEP="TRUE" *) reg [7:0] n457_q;
  (* KEEP="TRUE" *) wire n458_o;
  (* KEEP="TRUE" *) wire n459_o;
  (* KEEP="TRUE" *) wire n460_o;
  (* KEEP="TRUE" *) reg n461_q;
  (* KEEP="TRUE" *) wire [61:0] n462_o;
  (* KEEP="TRUE" *) wire [61:0] n463_o;
  (* KEEP="TRUE" *) wire [61:0] n464_o;
  (* KEEP="TRUE" *) reg [61:0] n465_q;
  (* KEEP="TRUE" *) wire [63:0] n467_o;
  (* KEEP="TRUE" *) reg [7:0] n468_q;
  (* KEEP="TRUE" *) reg [7:0] n469_q;
  (* KEEP="TRUE" *) reg [28:0] n470_q;
  (* KEEP="TRUE" *) wire [30:0] n471_o;
  (* KEEP="TRUE" *) reg [30:0] n472_q;
  (* KEEP="TRUE" *) wire [30:0] n473_o;
  (* KEEP="TRUE" *) reg [30:0] n474_q;
  (* KEEP="TRUE" *) reg [255:0] n475_q;
  (* KEEP="TRUE" *) reg [255:0] n476_q;
  (* KEEP="TRUE" *) reg n477_q;
  (* KEEP="TRUE" *) reg n478_q;
  (* KEEP="TRUE" *) reg n479_q;
  (* KEEP="TRUE" *) reg n480_q;
  (* KEEP="TRUE" *) wire n481_o;
  (* KEEP="TRUE" *) reg n482_q;
  (* KEEP="TRUE" *) reg [7:0] n483_q;
  (* KEEP="TRUE" *) reg [2:0] n484_q;
  (* KEEP="TRUE" *) wire [4:0] n485_o;
  (* KEEP="TRUE" *) reg [4:0] n486_q;
  (* KEEP="TRUE" *) reg n487_q;
  (* KEEP="TRUE" *) reg n488_q;
  (* KEEP="TRUE" *) reg n489_q;
  (* KEEP="TRUE" *) reg n490_q;
  (* KEEP="TRUE" *) reg n491_q;
  (* KEEP="TRUE" *) wire n493_data; // mem_rd
  (* KEEP="TRUE" *) wire n494_data; // mem_rd
  (* KEEP="TRUE" *) wire n495_data; // mem_rd
  (* KEEP="TRUE" *) wire n496_data; // mem_rd
  (* KEEP="TRUE" *) wire n497_o;
  (* KEEP="TRUE" *) wire n498_o;
  (* KEEP="TRUE" *) wire n499_o;
  (* KEEP="TRUE" *) wire n500_o;
  (* KEEP="TRUE" *) wire n501_o;
  (* KEEP="TRUE" *) wire n502_o;
  (* KEEP="TRUE" *) wire n503_o;
  (* KEEP="TRUE" *) wire n504_o;
  (* KEEP="TRUE" *) wire n505_o;
  (* KEEP="TRUE" *) wire n506_o;
  (* KEEP="TRUE" *) wire n507_o;
  (* KEEP="TRUE" *) wire n508_o;
  (* KEEP="TRUE" *) wire n509_o;
  (* KEEP="TRUE" *) wire n510_o;
  (* KEEP="TRUE" *) wire n511_o;
  (* KEEP="TRUE" *) wire n512_o;
  (* KEEP="TRUE" *) wire n513_o;
  (* KEEP="TRUE" *) wire n514_o;
  (* KEEP="TRUE" *) wire n515_o;
  (* KEEP="TRUE" *) wire n516_o;
  (* KEEP="TRUE" *) wire n517_o;
  (* KEEP="TRUE" *) wire n518_o;
  (* KEEP="TRUE" *) wire n519_o;
  (* KEEP="TRUE" *) wire n520_o;
  (* KEEP="TRUE" *) wire n521_o;
  (* KEEP="TRUE" *) wire n522_o;
  (* KEEP="TRUE" *) wire n523_o;
  (* KEEP="TRUE" *) wire n524_o;
  (* KEEP="TRUE" *) wire n525_o;
  (* KEEP="TRUE" *) wire n526_o;
  (* KEEP="TRUE" *) wire n527_o;
  (* KEEP="TRUE" *) wire n528_o;
  (* KEEP="TRUE" *) wire n529_o;
  (* KEEP="TRUE" *) wire n530_o;
  (* KEEP="TRUE" *) wire n531_o;
  (* KEEP="TRUE" *) wire n532_o;
  (* KEEP="TRUE" *) wire n533_o;
  (* KEEP="TRUE" *) wire n534_o;
  (* KEEP="TRUE" *) wire n535_o;
  (* KEEP="TRUE" *) wire n536_o;
  (* KEEP="TRUE" *) wire n537_o;
  (* KEEP="TRUE" *) wire n538_o;
  (* KEEP="TRUE" *) wire n539_o;
  (* KEEP="TRUE" *) wire n540_o;
  (* KEEP="TRUE" *) wire n541_o;
  (* KEEP="TRUE" *) wire n542_o;
  (* KEEP="TRUE" *) wire n543_o;
  (* KEEP="TRUE" *) wire n544_o;
  (* KEEP="TRUE" *) wire n545_o;
  (* KEEP="TRUE" *) wire n546_o;
  (* KEEP="TRUE" *) wire n547_o;
  (* KEEP="TRUE" *) wire n548_o;
  (* KEEP="TRUE" *) wire n549_o;
  (* KEEP="TRUE" *) wire n550_o;
  (* KEEP="TRUE" *) wire n551_o;
  (* KEEP="TRUE" *) wire n552_o;
  (* KEEP="TRUE" *) wire n553_o;
  (* KEEP="TRUE" *) wire n554_o;
  (* KEEP="TRUE" *) wire n555_o;
  (* KEEP="TRUE" *) wire n556_o;
  (* KEEP="TRUE" *) wire n557_o;
  (* KEEP="TRUE" *) wire n558_o;
  (* KEEP="TRUE" *) wire n559_o;
  (* KEEP="TRUE" *) wire n560_o;
  (* KEEP="TRUE" *) wire n561_o;
  (* KEEP="TRUE" *) wire n562_o;
  (* KEEP="TRUE" *) wire n563_o;
  (* KEEP="TRUE" *) wire n564_o;
  (* KEEP="TRUE" *) wire n565_o;
  (* KEEP="TRUE" *) wire n566_o;
  (* KEEP="TRUE" *) wire n567_o;
  (* KEEP="TRUE" *) wire n568_o;
  (* KEEP="TRUE" *) wire n569_o;
  (* KEEP="TRUE" *) wire n570_o;
  (* KEEP="TRUE" *) wire n571_o;
  (* KEEP="TRUE" *) wire n572_o;
  (* KEEP="TRUE" *) wire n573_o;
  (* KEEP="TRUE" *) wire n574_o;
  (* KEEP="TRUE" *) wire n575_o;
  (* KEEP="TRUE" *) wire n576_o;
  (* KEEP="TRUE" *) wire n577_o;
  (* KEEP="TRUE" *) wire n578_o;
  (* KEEP="TRUE" *) wire n579_o;
  (* KEEP="TRUE" *) wire n580_o;
  (* KEEP="TRUE" *) wire n581_o;
  (* KEEP="TRUE" *) wire n582_o;
  (* KEEP="TRUE" *) wire n583_o;
  (* KEEP="TRUE" *) wire n584_o;
  (* KEEP="TRUE" *) wire n585_o;
  (* KEEP="TRUE" *) wire n586_o;
  (* KEEP="TRUE" *) wire n587_o;
  (* KEEP="TRUE" *) wire n588_o;
  (* KEEP="TRUE" *) wire n589_o;
  (* KEEP="TRUE" *) wire n590_o;
  (* KEEP="TRUE" *) wire n591_o;
  (* KEEP="TRUE" *) wire n592_o;
  (* KEEP="TRUE" *) wire n593_o;
  (* KEEP="TRUE" *) wire n594_o;
  (* KEEP="TRUE" *) wire n595_o;
  (* KEEP="TRUE" *) wire n596_o;
  (* KEEP="TRUE" *) wire n597_o;
  (* KEEP="TRUE" *) wire n598_o;
  (* KEEP="TRUE" *) wire n599_o;
  (* KEEP="TRUE" *) wire n600_o;
  (* KEEP="TRUE" *) wire n601_o;
  (* KEEP="TRUE" *) wire n602_o;
  (* KEEP="TRUE" *) wire n603_o;
  (* KEEP="TRUE" *) wire n604_o;
  (* KEEP="TRUE" *) wire n605_o;
  (* KEEP="TRUE" *) wire n606_o;
  (* KEEP="TRUE" *) wire n607_o;
  (* KEEP="TRUE" *) wire n608_o;
  (* KEEP="TRUE" *) wire n609_o;
  (* KEEP="TRUE" *) wire n610_o;
  (* KEEP="TRUE" *) wire n611_o;
  (* KEEP="TRUE" *) wire n612_o;
  (* KEEP="TRUE" *) wire n613_o;
  (* KEEP="TRUE" *) wire n614_o;
  (* KEEP="TRUE" *) wire n615_o;
  (* KEEP="TRUE" *) wire n616_o;
  (* KEEP="TRUE" *) wire n617_o;
  (* KEEP="TRUE" *) wire n618_o;
  (* KEEP="TRUE" *) wire n619_o;
  (* KEEP="TRUE" *) wire n620_o;
  (* KEEP="TRUE" *) wire n621_o;
  (* KEEP="TRUE" *) wire n622_o;
  (* KEEP="TRUE" *) wire n623_o;
  (* KEEP="TRUE" *) wire n624_o;
  (* KEEP="TRUE" *) wire n625_o;
  (* KEEP="TRUE" *) wire n626_o;
  (* KEEP="TRUE" *) wire n627_o;
  (* KEEP="TRUE" *) wire n628_o;
  (* KEEP="TRUE" *) wire n629_o;
  (* KEEP="TRUE" *) wire n630_o;
  (* KEEP="TRUE" *) wire n631_o;
  (* KEEP="TRUE" *) wire n632_o;
  (* KEEP="TRUE" *) wire n633_o;
  (* KEEP="TRUE" *) wire n634_o;
  (* KEEP="TRUE" *) wire n635_o;
  (* KEEP="TRUE" *) wire n636_o;
  (* KEEP="TRUE" *) wire n637_o;
  (* KEEP="TRUE" *) wire n638_o;
  (* KEEP="TRUE" *) wire n639_o;
  (* KEEP="TRUE" *) wire n640_o;
  (* KEEP="TRUE" *) wire n641_o;
  (* KEEP="TRUE" *) wire n642_o;
  (* KEEP="TRUE" *) wire n643_o;
  (* KEEP="TRUE" *) wire n644_o;
  (* KEEP="TRUE" *) wire n645_o;
  (* KEEP="TRUE" *) wire n646_o;
  (* KEEP="TRUE" *) wire n647_o;
  (* KEEP="TRUE" *) wire n648_o;
  (* KEEP="TRUE" *) wire n649_o;
  (* KEEP="TRUE" *) wire n650_o;
  (* KEEP="TRUE" *) wire n651_o;
  (* KEEP="TRUE" *) wire n652_o;
  (* KEEP="TRUE" *) wire n653_o;
  (* KEEP="TRUE" *) wire n654_o;
  (* KEEP="TRUE" *) wire n655_o;
  (* KEEP="TRUE" *) wire n656_o;
  (* KEEP="TRUE" *) wire n657_o;
  (* KEEP="TRUE" *) wire n658_o;
  (* KEEP="TRUE" *) wire n659_o;
  (* KEEP="TRUE" *) wire n660_o;
  (* KEEP="TRUE" *) wire n661_o;
  (* KEEP="TRUE" *) wire n662_o;
  (* KEEP="TRUE" *) wire n663_o;
  (* KEEP="TRUE" *) wire n664_o;
  (* KEEP="TRUE" *) wire n665_o;
  (* KEEP="TRUE" *) wire n666_o;
  (* KEEP="TRUE" *) wire n667_o;
  (* KEEP="TRUE" *) wire n668_o;
  (* KEEP="TRUE" *) wire n669_o;
  (* KEEP="TRUE" *) wire n670_o;
  (* KEEP="TRUE" *) wire n671_o;
  (* KEEP="TRUE" *) wire n672_o;
  (* KEEP="TRUE" *) wire n673_o;
  (* KEEP="TRUE" *) wire n674_o;
  (* KEEP="TRUE" *) wire n675_o;
  (* KEEP="TRUE" *) wire n676_o;
  (* KEEP="TRUE" *) wire n677_o;
  (* KEEP="TRUE" *) wire n678_o;
  (* KEEP="TRUE" *) wire n679_o;
  (* KEEP="TRUE" *) wire n680_o;
  (* KEEP="TRUE" *) wire n681_o;
  (* KEEP="TRUE" *) wire n682_o;
  (* KEEP="TRUE" *) wire n683_o;
  (* KEEP="TRUE" *) wire n684_o;
  (* KEEP="TRUE" *) wire n685_o;
  (* KEEP="TRUE" *) wire n686_o;
  (* KEEP="TRUE" *) wire n687_o;
  (* KEEP="TRUE" *) wire n688_o;
  (* KEEP="TRUE" *) wire n689_o;
  (* KEEP="TRUE" *) wire n690_o;
  (* KEEP="TRUE" *) wire n691_o;
  (* KEEP="TRUE" *) wire n692_o;
  (* KEEP="TRUE" *) wire n693_o;
  (* KEEP="TRUE" *) wire n694_o;
  (* KEEP="TRUE" *) wire n695_o;
  (* KEEP="TRUE" *) wire n696_o;
  (* KEEP="TRUE" *) wire n697_o;
  (* KEEP="TRUE" *) wire n698_o;
  (* KEEP="TRUE" *) wire n699_o;
  (* KEEP="TRUE" *) wire n700_o;
  (* KEEP="TRUE" *) wire n701_o;
  (* KEEP="TRUE" *) wire n702_o;
  (* KEEP="TRUE" *) wire n703_o;
  (* KEEP="TRUE" *) wire n704_o;
  (* KEEP="TRUE" *) wire n705_o;
  (* KEEP="TRUE" *) wire n706_o;
  (* KEEP="TRUE" *) wire n707_o;
  (* KEEP="TRUE" *) wire n708_o;
  (* KEEP="TRUE" *) wire n709_o;
  (* KEEP="TRUE" *) wire n710_o;
  (* KEEP="TRUE" *) wire n711_o;
  (* KEEP="TRUE" *) wire n712_o;
  (* KEEP="TRUE" *) wire n713_o;
  (* KEEP="TRUE" *) wire n714_o;
  (* KEEP="TRUE" *) wire n715_o;
  (* KEEP="TRUE" *) wire n716_o;
  (* KEEP="TRUE" *) wire n717_o;
  (* KEEP="TRUE" *) wire n718_o;
  (* KEEP="TRUE" *) wire n719_o;
  (* KEEP="TRUE" *) wire n720_o;
  (* KEEP="TRUE" *) wire n721_o;
  (* KEEP="TRUE" *) wire n722_o;
  (* KEEP="TRUE" *) wire n723_o;
  (* KEEP="TRUE" *) wire n724_o;
  (* KEEP="TRUE" *) wire n725_o;
  (* KEEP="TRUE" *) wire n726_o;
  (* KEEP="TRUE" *) wire n727_o;
  (* KEEP="TRUE" *) wire n728_o;
  (* KEEP="TRUE" *) wire n729_o;
  (* KEEP="TRUE" *) wire n730_o;
  (* KEEP="TRUE" *) wire n731_o;
  (* KEEP="TRUE" *) wire n732_o;
  (* KEEP="TRUE" *) wire n733_o;
  (* KEEP="TRUE" *) wire n734_o;
  (* KEEP="TRUE" *) wire n735_o;
  (* KEEP="TRUE" *) wire n736_o;
  (* KEEP="TRUE" *) wire n737_o;
  (* KEEP="TRUE" *) wire n738_o;
  (* KEEP="TRUE" *) wire n739_o;
  (* KEEP="TRUE" *) wire n740_o;
  (* KEEP="TRUE" *) wire n741_o;
  (* KEEP="TRUE" *) wire n742_o;
  (* KEEP="TRUE" *) wire n743_o;
  (* KEEP="TRUE" *) wire n744_o;
  (* KEEP="TRUE" *) wire n745_o;
  (* KEEP="TRUE" *) wire n746_o;
  (* KEEP="TRUE" *) wire n747_o;
  (* KEEP="TRUE" *) wire n748_o;
  (* KEEP="TRUE" *) wire n749_o;
  (* KEEP="TRUE" *) wire n750_o;
  (* KEEP="TRUE" *) wire n751_o;
  (* KEEP="TRUE" *) wire n752_o;
  (* KEEP="TRUE" *) wire n753_o;
  (* KEEP="TRUE" *) wire n754_o;
  (* KEEP="TRUE" *) wire n755_o;
  (* KEEP="TRUE" *) wire n756_o;
  (* KEEP="TRUE" *) wire n757_o;
  (* KEEP="TRUE" *) wire n758_o;
  (* KEEP="TRUE" *) wire n759_o;
  (* KEEP="TRUE" *) wire n760_o;
  (* KEEP="TRUE" *) wire n761_o;
  (* KEEP="TRUE" *) wire n762_o;
  (* KEEP="TRUE" *) wire n763_o;
  (* KEEP="TRUE" *) wire n764_o;
  (* KEEP="TRUE" *) wire n765_o;
  (* KEEP="TRUE" *) wire n766_o;
  (* KEEP="TRUE" *) wire n767_o;
  (* KEEP="TRUE" *) wire n768_o;
  (* KEEP="TRUE" *) wire n769_o;
  (* KEEP="TRUE" *) wire n770_o;
  (* KEEP="TRUE" *) wire n771_o;
  (* KEEP="TRUE" *) wire n772_o;
  (* KEEP="TRUE" *) wire n773_o;
  (* KEEP="TRUE" *) wire n774_o;
  (* KEEP="TRUE" *) wire n775_o;
  (* KEEP="TRUE" *) wire n776_o;
  (* KEEP="TRUE" *) wire n777_o;
  (* KEEP="TRUE" *) wire n778_o;
  (* KEEP="TRUE" *) wire n779_o;
  (* KEEP="TRUE" *) wire n780_o;
  (* KEEP="TRUE" *) wire n781_o;
  (* KEEP="TRUE" *) wire n782_o;
  (* KEEP="TRUE" *) wire n783_o;
  (* KEEP="TRUE" *) wire n784_o;
  (* KEEP="TRUE" *) wire n785_o;
  (* KEEP="TRUE" *) wire n786_o;
  (* KEEP="TRUE" *) wire n787_o;
  (* KEEP="TRUE" *) wire n788_o;
  (* KEEP="TRUE" *) wire n789_o;
  (* KEEP="TRUE" *) wire n790_o;
  (* KEEP="TRUE" *) wire n791_o;
  (* KEEP="TRUE" *) wire n792_o;
  (* KEEP="TRUE" *) wire n793_o;
  (* KEEP="TRUE" *) wire n794_o;
  (* KEEP="TRUE" *) wire n795_o;
  (* KEEP="TRUE" *) wire n796_o;
  (* KEEP="TRUE" *) wire n797_o;
  (* KEEP="TRUE" *) wire n798_o;
  (* KEEP="TRUE" *) wire n799_o;
  (* KEEP="TRUE" *) wire n800_o;
  (* KEEP="TRUE" *) wire n801_o;
  (* KEEP="TRUE" *) wire n802_o;
  (* KEEP="TRUE" *) wire n803_o;
  (* KEEP="TRUE" *) wire n804_o;
  (* KEEP="TRUE" *) wire n805_o;
  (* KEEP="TRUE" *) wire n806_o;
  (* KEEP="TRUE" *) wire n807_o;
  (* KEEP="TRUE" *) wire n808_o;
  (* KEEP="TRUE" *) wire n809_o;
  (* KEEP="TRUE" *) wire n810_o;
  (* KEEP="TRUE" *) wire n811_o;
  (* KEEP="TRUE" *) wire n812_o;
  (* KEEP="TRUE" *) wire n813_o;
  (* KEEP="TRUE" *) wire n814_o;
  (* KEEP="TRUE" *) wire n815_o;
  (* KEEP="TRUE" *) wire n816_o;
  (* KEEP="TRUE" *) wire n817_o;
  (* KEEP="TRUE" *) wire n818_o;
  (* KEEP="TRUE" *) wire n819_o;
  (* KEEP="TRUE" *) wire n820_o;
  (* KEEP="TRUE" *) wire n821_o;
  (* KEEP="TRUE" *) wire n822_o;
  (* KEEP="TRUE" *) wire n823_o;
  (* KEEP="TRUE" *) wire n824_o;
  (* KEEP="TRUE" *) wire n825_o;
  (* KEEP="TRUE" *) wire n826_o;
  (* KEEP="TRUE" *) wire n827_o;
  (* KEEP="TRUE" *) wire n828_o;
  (* KEEP="TRUE" *) wire n829_o;
  (* KEEP="TRUE" *) wire n830_o;
  (* KEEP="TRUE" *) wire n831_o;
  (* KEEP="TRUE" *) wire n832_o;
  (* KEEP="TRUE" *) wire n833_o;
  (* KEEP="TRUE" *) wire n834_o;
  (* KEEP="TRUE" *) wire n835_o;
  (* KEEP="TRUE" *) wire n836_o;
  (* KEEP="TRUE" *) wire n837_o;
  (* KEEP="TRUE" *) wire n838_o;
  (* KEEP="TRUE" *) wire n839_o;
  (* KEEP="TRUE" *) wire n840_o;
  (* KEEP="TRUE" *) wire n841_o;
  (* KEEP="TRUE" *) wire n842_o;
  (* KEEP="TRUE" *) wire n843_o;
  (* KEEP="TRUE" *) wire n844_o;
  (* KEEP="TRUE" *) wire n845_o;
  (* KEEP="TRUE" *) wire n846_o;
  (* KEEP="TRUE" *) wire n847_o;
  (* KEEP="TRUE" *) wire n848_o;
  (* KEEP="TRUE" *) wire n849_o;
  (* KEEP="TRUE" *) wire n850_o;
  (* KEEP="TRUE" *) wire n851_o;
  (* KEEP="TRUE" *) wire n852_o;
  (* KEEP="TRUE" *) wire n853_o;
  (* KEEP="TRUE" *) wire n854_o;
  (* KEEP="TRUE" *) wire n855_o;
  (* KEEP="TRUE" *) wire n856_o;
  (* KEEP="TRUE" *) wire n857_o;
  (* KEEP="TRUE" *) wire n858_o;
  (* KEEP="TRUE" *) wire n859_o;
  (* KEEP="TRUE" *) wire n860_o;
  (* KEEP="TRUE" *) wire n861_o;
  (* KEEP="TRUE" *) wire n862_o;
  (* KEEP="TRUE" *) wire n863_o;
  (* KEEP="TRUE" *) wire n864_o;
  (* KEEP="TRUE" *) wire n865_o;
  (* KEEP="TRUE" *) wire n866_o;
  (* KEEP="TRUE" *) wire n867_o;
  (* KEEP="TRUE" *) wire n868_o;
  (* KEEP="TRUE" *) wire n869_o;
  (* KEEP="TRUE" *) wire n870_o;
  (* KEEP="TRUE" *) wire n871_o;
  (* KEEP="TRUE" *) wire n872_o;
  (* KEEP="TRUE" *) wire n873_o;
  (* KEEP="TRUE" *) wire n874_o;
  (* KEEP="TRUE" *) wire n875_o;
  (* KEEP="TRUE" *) wire n876_o;
  (* KEEP="TRUE" *) wire n877_o;
  (* KEEP="TRUE" *) wire n878_o;
  (* KEEP="TRUE" *) wire n879_o;
  (* KEEP="TRUE" *) wire n880_o;
  (* KEEP="TRUE" *) wire n881_o;
  (* KEEP="TRUE" *) wire n882_o;
  (* KEEP="TRUE" *) wire n883_o;
  (* KEEP="TRUE" *) wire n884_o;
  (* KEEP="TRUE" *) wire n885_o;
  (* KEEP="TRUE" *) wire n886_o;
  (* KEEP="TRUE" *) wire n887_o;
  (* KEEP="TRUE" *) wire n888_o;
  (* KEEP="TRUE" *) wire n889_o;
  (* KEEP="TRUE" *) wire n890_o;
  (* KEEP="TRUE" *) wire n891_o;
  (* KEEP="TRUE" *) wire n892_o;
  (* KEEP="TRUE" *) wire n893_o;
  (* KEEP="TRUE" *) wire n894_o;
  (* KEEP="TRUE" *) wire n895_o;
  (* KEEP="TRUE" *) wire n896_o;
  (* KEEP="TRUE" *) wire n897_o;
  (* KEEP="TRUE" *) wire n898_o;
  (* KEEP="TRUE" *) wire n899_o;
  (* KEEP="TRUE" *) wire n900_o;
  (* KEEP="TRUE" *) wire n901_o;
  (* KEEP="TRUE" *) wire n902_o;
  (* KEEP="TRUE" *) wire n903_o;
  (* KEEP="TRUE" *) wire n904_o;
  (* KEEP="TRUE" *) wire n905_o;
  (* KEEP="TRUE" *) wire n906_o;
  (* KEEP="TRUE" *) wire n907_o;
  (* KEEP="TRUE" *) wire n908_o;
  (* KEEP="TRUE" *) wire n909_o;
  (* KEEP="TRUE" *) wire n910_o;
  (* KEEP="TRUE" *) wire n911_o;
  (* KEEP="TRUE" *) wire n912_o;
  (* KEEP="TRUE" *) wire n913_o;
  (* KEEP="TRUE" *) wire n914_o;
  (* KEEP="TRUE" *) wire n915_o;
  (* KEEP="TRUE" *) wire n916_o;
  (* KEEP="TRUE" *) wire n917_o;
  (* KEEP="TRUE" *) wire n918_o;
  (* KEEP="TRUE" *) wire n919_o;
  (* KEEP="TRUE" *) wire n920_o;
  (* KEEP="TRUE" *) wire n921_o;
  (* KEEP="TRUE" *) wire n922_o;
  (* KEEP="TRUE" *) wire n923_o;
  (* KEEP="TRUE" *) wire n924_o;
  (* KEEP="TRUE" *) wire n925_o;
  (* KEEP="TRUE" *) wire n926_o;
  (* KEEP="TRUE" *) wire n927_o;
  (* KEEP="TRUE" *) wire n928_o;
  (* KEEP="TRUE" *) wire n929_o;
  (* KEEP="TRUE" *) wire n930_o;
  (* KEEP="TRUE" *) wire n931_o;
  (* KEEP="TRUE" *) wire n932_o;
  (* KEEP="TRUE" *) wire n933_o;
  (* KEEP="TRUE" *) wire n934_o;
  (* KEEP="TRUE" *) wire n935_o;
  (* KEEP="TRUE" *) wire n936_o;
  (* KEEP="TRUE" *) wire n937_o;
  (* KEEP="TRUE" *) wire n938_o;
  (* KEEP="TRUE" *) wire n939_o;
  (* KEEP="TRUE" *) wire n940_o;
  (* KEEP="TRUE" *) wire n941_o;
  (* KEEP="TRUE" *) wire n942_o;
  (* KEEP="TRUE" *) wire n943_o;
  (* KEEP="TRUE" *) wire n944_o;
  (* KEEP="TRUE" *) wire n945_o;
  (* KEEP="TRUE" *) wire n946_o;
  (* KEEP="TRUE" *) wire n947_o;
  (* KEEP="TRUE" *) wire n948_o;
  (* KEEP="TRUE" *) wire n949_o;
  (* KEEP="TRUE" *) wire n950_o;
  (* KEEP="TRUE" *) wire n951_o;
  (* KEEP="TRUE" *) wire n952_o;
  (* KEEP="TRUE" *) wire n953_o;
  (* KEEP="TRUE" *) wire n954_o;
  (* KEEP="TRUE" *) wire n955_o;
  (* KEEP="TRUE" *) wire n956_o;
  (* KEEP="TRUE" *) wire n957_o;
  (* KEEP="TRUE" *) wire n958_o;
  (* KEEP="TRUE" *) wire n959_o;
  (* KEEP="TRUE" *) wire n960_o;
  (* KEEP="TRUE" *) wire n961_o;
  (* KEEP="TRUE" *) wire n962_o;
  (* KEEP="TRUE" *) wire n963_o;
  (* KEEP="TRUE" *) wire n964_o;
  (* KEEP="TRUE" *) wire n965_o;
  (* KEEP="TRUE" *) wire n966_o;
  (* KEEP="TRUE" *) wire n967_o;
  (* KEEP="TRUE" *) wire n968_o;
  (* KEEP="TRUE" *) wire n969_o;
  (* KEEP="TRUE" *) wire n970_o;
  (* KEEP="TRUE" *) wire n971_o;
  (* KEEP="TRUE" *) wire n972_o;
  (* KEEP="TRUE" *) wire n973_o;
  (* KEEP="TRUE" *) wire n974_o;
  (* KEEP="TRUE" *) wire n975_o;
  (* KEEP="TRUE" *) wire n976_o;
  (* KEEP="TRUE" *) wire n977_o;
  (* KEEP="TRUE" *) wire n978_o;
  (* KEEP="TRUE" *) wire n979_o;
  (* KEEP="TRUE" *) wire n980_o;
  (* KEEP="TRUE" *) wire n981_o;
  (* KEEP="TRUE" *) wire n982_o;
  (* KEEP="TRUE" *) wire n983_o;
  (* KEEP="TRUE" *) wire n984_o;
  (* KEEP="TRUE" *) wire n985_o;
  (* KEEP="TRUE" *) wire n986_o;
  (* KEEP="TRUE" *) wire n987_o;
  (* KEEP="TRUE" *) wire n988_o;
  (* KEEP="TRUE" *) wire n989_o;
  (* KEEP="TRUE" *) wire n990_o;
  (* KEEP="TRUE" *) wire n991_o;
  (* KEEP="TRUE" *) wire n992_o;
  (* KEEP="TRUE" *) wire n993_o;
  (* KEEP="TRUE" *) wire n994_o;
  (* KEEP="TRUE" *) wire n995_o;
  (* KEEP="TRUE" *) wire n996_o;
  (* KEEP="TRUE" *) wire n997_o;
  (* KEEP="TRUE" *) wire n998_o;
  (* KEEP="TRUE" *) wire n999_o;
  (* KEEP="TRUE" *) wire n1000_o;
  (* KEEP="TRUE" *) wire n1001_o;
  (* KEEP="TRUE" *) wire n1002_o;
  (* KEEP="TRUE" *) wire n1003_o;
  (* KEEP="TRUE" *) wire n1004_o;
  (* KEEP="TRUE" *) wire n1005_o;
  (* KEEP="TRUE" *) wire n1006_o;
  (* KEEP="TRUE" *) wire n1007_o;
  (* KEEP="TRUE" *) wire n1008_o;
  (* KEEP="TRUE" *) wire n1009_o;
  (* KEEP="TRUE" *) wire n1010_o;
  (* KEEP="TRUE" *) wire n1011_o;
  (* KEEP="TRUE" *) wire n1012_o;
  (* KEEP="TRUE" *) wire n1013_o;
  (* KEEP="TRUE" *) wire n1014_o;
  (* KEEP="TRUE" *) wire n1015_o;
  (* KEEP="TRUE" *) wire n1016_o;
  (* KEEP="TRUE" *) wire n1017_o;
  (* KEEP="TRUE" *) wire n1018_o;
  (* KEEP="TRUE" *) wire n1019_o;
  (* KEEP="TRUE" *) wire n1020_o;
  (* KEEP="TRUE" *) wire n1021_o;
  (* KEEP="TRUE" *) wire n1022_o;
  (* KEEP="TRUE" *) wire n1023_o;
  (* KEEP="TRUE" *) wire n1024_o;
  (* KEEP="TRUE" *) wire n1025_o;
  (* KEEP="TRUE" *) wire n1026_o;
  (* KEEP="TRUE" *) wire n1027_o;
  (* KEEP="TRUE" *) wire n1028_o;
  (* KEEP="TRUE" *) wire n1029_o;
  (* KEEP="TRUE" *) wire n1030_o;
  (* KEEP="TRUE" *) wire n1031_o;
  (* KEEP="TRUE" *) wire n1032_o;
  (* KEEP="TRUE" *) wire n1033_o;
  (* KEEP="TRUE" *) wire n1034_o;
  (* KEEP="TRUE" *) wire n1035_o;
  (* KEEP="TRUE" *) wire n1036_o;
  (* KEEP="TRUE" *) wire n1037_o;
  (* KEEP="TRUE" *) wire n1038_o;
  (* KEEP="TRUE" *) wire n1039_o;
  (* KEEP="TRUE" *) wire n1040_o;
  (* KEEP="TRUE" *) wire n1041_o;
  (* KEEP="TRUE" *) wire n1042_o;
  (* KEEP="TRUE" *) wire n1043_o;
  (* KEEP="TRUE" *) wire n1044_o;
  (* KEEP="TRUE" *) wire n1045_o;
  (* KEEP="TRUE" *) wire n1046_o;
  (* KEEP="TRUE" *) wire n1047_o;
  (* KEEP="TRUE" *) wire n1048_o;
  (* KEEP="TRUE" *) wire n1049_o;
  (* KEEP="TRUE" *) wire n1050_o;
  (* KEEP="TRUE" *) wire n1051_o;
  (* KEEP="TRUE" *) wire n1052_o;
  (* KEEP="TRUE" *) wire n1053_o;
  (* KEEP="TRUE" *) wire n1054_o;
  (* KEEP="TRUE" *) wire n1055_o;
  (* KEEP="TRUE" *) wire n1056_o;
  (* KEEP="TRUE" *) wire n1057_o;
  (* KEEP="TRUE" *) wire n1058_o;
  (* KEEP="TRUE" *) wire n1059_o;
  (* KEEP="TRUE" *) wire n1060_o;
  (* KEEP="TRUE" *) wire n1061_o;
  (* KEEP="TRUE" *) wire n1062_o;
  (* KEEP="TRUE" *) wire n1063_o;
  (* KEEP="TRUE" *) wire n1064_o;
  (* KEEP="TRUE" *) wire n1065_o;
  (* KEEP="TRUE" *) wire n1066_o;
  (* KEEP="TRUE" *) wire n1067_o;
  (* KEEP="TRUE" *) wire n1068_o;
  (* KEEP="TRUE" *) wire n1069_o;
  (* KEEP="TRUE" *) wire n1070_o;
  (* KEEP="TRUE" *) wire n1071_o;
  (* KEEP="TRUE" *) wire n1072_o;
  (* KEEP="TRUE" *) wire n1073_o;
  (* KEEP="TRUE" *) wire n1074_o;
  (* KEEP="TRUE" *) wire n1075_o;
  (* KEEP="TRUE" *) wire n1076_o;
  (* KEEP="TRUE" *) wire n1077_o;
  (* KEEP="TRUE" *) wire n1078_o;
  (* KEEP="TRUE" *) wire n1079_o;
  (* KEEP="TRUE" *) wire n1080_o;
  (* KEEP="TRUE" *) wire n1081_o;
  (* KEEP="TRUE" *) wire n1082_o;
  (* KEEP="TRUE" *) wire n1083_o;
  (* KEEP="TRUE" *) wire n1084_o;
  (* KEEP="TRUE" *) wire n1085_o;
  (* KEEP="TRUE" *) wire n1086_o;
  (* KEEP="TRUE" *) wire n1087_o;
  (* KEEP="TRUE" *) wire n1088_o;
  (* KEEP="TRUE" *) wire n1089_o;
  (* KEEP="TRUE" *) wire n1090_o;
  (* KEEP="TRUE" *) wire n1091_o;
  (* KEEP="TRUE" *) wire n1092_o;
  (* KEEP="TRUE" *) wire n1093_o;
  (* KEEP="TRUE" *) wire n1094_o;
  (* KEEP="TRUE" *) wire n1095_o;
  (* KEEP="TRUE" *) wire n1096_o;
  (* KEEP="TRUE" *) wire n1097_o;
  (* KEEP="TRUE" *) wire n1098_o;
  (* KEEP="TRUE" *) wire n1099_o;
  (* KEEP="TRUE" *) wire n1100_o;
  (* KEEP="TRUE" *) wire n1101_o;
  (* KEEP="TRUE" *) wire n1102_o;
  (* KEEP="TRUE" *) wire n1103_o;
  (* KEEP="TRUE" *) wire n1104_o;
  (* KEEP="TRUE" *) wire n1105_o;
  (* KEEP="TRUE" *) wire n1106_o;
  (* KEEP="TRUE" *) wire n1107_o;
  (* KEEP="TRUE" *) wire n1108_o;
  (* KEEP="TRUE" *) wire n1109_o;
  (* KEEP="TRUE" *) wire n1110_o;
  (* KEEP="TRUE" *) wire n1111_o;
  (* KEEP="TRUE" *) wire n1112_o;
  (* KEEP="TRUE" *) wire n1113_o;
  (* KEEP="TRUE" *) wire n1114_o;
  (* KEEP="TRUE" *) wire n1115_o;
  (* KEEP="TRUE" *) wire n1116_o;
  (* KEEP="TRUE" *) wire n1117_o;
  (* KEEP="TRUE" *) wire n1118_o;
  (* KEEP="TRUE" *) wire n1119_o;
  (* KEEP="TRUE" *) wire n1120_o;
  (* KEEP="TRUE" *) wire n1121_o;
  (* KEEP="TRUE" *) wire n1122_o;
  (* KEEP="TRUE" *) wire n1123_o;
  (* KEEP="TRUE" *) wire n1124_o;
  (* KEEP="TRUE" *) wire n1125_o;
  (* KEEP="TRUE" *) wire n1126_o;
  (* KEEP="TRUE" *) wire n1127_o;
  (* KEEP="TRUE" *) wire n1128_o;
  (* KEEP="TRUE" *) wire n1129_o;
  (* KEEP="TRUE" *) wire n1130_o;
  (* KEEP="TRUE" *) wire n1131_o;
  (* KEEP="TRUE" *) wire n1132_o;
  (* KEEP="TRUE" *) wire n1133_o;
  (* KEEP="TRUE" *) wire n1134_o;
  (* KEEP="TRUE" *) wire n1135_o;
  (* KEEP="TRUE" *) wire n1136_o;
  (* KEEP="TRUE" *) wire n1137_o;
  (* KEEP="TRUE" *) wire n1138_o;
  (* KEEP="TRUE" *) wire n1139_o;
  (* KEEP="TRUE" *) wire n1140_o;
  (* KEEP="TRUE" *) wire n1141_o;
  (* KEEP="TRUE" *) wire n1142_o;
  (* KEEP="TRUE" *) wire n1143_o;
  (* KEEP="TRUE" *) wire n1144_o;
  (* KEEP="TRUE" *) wire n1145_o;
  (* KEEP="TRUE" *) wire n1146_o;
  (* KEEP="TRUE" *) wire n1147_o;
  (* KEEP="TRUE" *) wire n1148_o;
  (* KEEP="TRUE" *) wire n1149_o;
  (* KEEP="TRUE" *) wire n1150_o;
  (* KEEP="TRUE" *) wire n1151_o;
  (* KEEP="TRUE" *) wire n1152_o;
  (* KEEP="TRUE" *) wire n1153_o;
  (* KEEP="TRUE" *) wire n1154_o;
  (* KEEP="TRUE" *) wire n1155_o;
  (* KEEP="TRUE" *) wire n1156_o;
  (* KEEP="TRUE" *) wire n1157_o;
  (* KEEP="TRUE" *) wire n1158_o;
  (* KEEP="TRUE" *) wire n1159_o;
  (* KEEP="TRUE" *) wire n1160_o;
  (* KEEP="TRUE" *) wire n1161_o;
  (* KEEP="TRUE" *) wire n1162_o;
  (* KEEP="TRUE" *) wire n1163_o;
  (* KEEP="TRUE" *) wire n1164_o;
  (* KEEP="TRUE" *) wire n1165_o;
  (* KEEP="TRUE" *) wire n1166_o;
  (* KEEP="TRUE" *) wire n1167_o;
  (* KEEP="TRUE" *) wire n1168_o;
  (* KEEP="TRUE" *) wire n1169_o;
  (* KEEP="TRUE" *) wire n1170_o;
  (* KEEP="TRUE" *) wire n1171_o;
  (* KEEP="TRUE" *) wire n1172_o;
  (* KEEP="TRUE" *) wire n1173_o;
  (* KEEP="TRUE" *) wire n1174_o;
  (* KEEP="TRUE" *) wire n1175_o;
  (* KEEP="TRUE" *) wire n1176_o;
  (* KEEP="TRUE" *) wire n1177_o;
  (* KEEP="TRUE" *) wire n1178_o;
  (* KEEP="TRUE" *) wire n1179_o;
  (* KEEP="TRUE" *) wire n1180_o;
  (* KEEP="TRUE" *) wire n1181_o;
  (* KEEP="TRUE" *) wire n1182_o;
  (* KEEP="TRUE" *) wire n1183_o;
  (* KEEP="TRUE" *) wire n1184_o;
  (* KEEP="TRUE" *) wire n1185_o;
  (* KEEP="TRUE" *) wire n1186_o;
  (* KEEP="TRUE" *) wire n1187_o;
  (* KEEP="TRUE" *) wire n1188_o;
  (* KEEP="TRUE" *) wire n1189_o;
  (* KEEP="TRUE" *) wire n1190_o;
  (* KEEP="TRUE" *) wire n1191_o;
  (* KEEP="TRUE" *) wire n1192_o;
  (* KEEP="TRUE" *) wire n1193_o;
  (* KEEP="TRUE" *) wire n1194_o;
  (* KEEP="TRUE" *) wire n1195_o;
  (* KEEP="TRUE" *) wire n1196_o;
  (* KEEP="TRUE" *) wire n1197_o;
  (* KEEP="TRUE" *) wire n1198_o;
  (* KEEP="TRUE" *) wire n1199_o;
  (* KEEP="TRUE" *) wire n1200_o;
  (* KEEP="TRUE" *) wire n1201_o;
  (* KEEP="TRUE" *) wire n1202_o;
  (* KEEP="TRUE" *) wire n1203_o;
  (* KEEP="TRUE" *) wire n1204_o;
  (* KEEP="TRUE" *) wire n1205_o;
  (* KEEP="TRUE" *) wire n1206_o;
  (* KEEP="TRUE" *) wire n1207_o;
  (* KEEP="TRUE" *) wire n1208_o;
  (* KEEP="TRUE" *) wire n1209_o;
  (* KEEP="TRUE" *) wire n1210_o;
  (* KEEP="TRUE" *) wire n1211_o;
  (* KEEP="TRUE" *) wire n1212_o;
  (* KEEP="TRUE" *) wire n1213_o;
  (* KEEP="TRUE" *) wire n1214_o;
  (* KEEP="TRUE" *) wire n1215_o;
  (* KEEP="TRUE" *) wire n1216_o;
  (* KEEP="TRUE" *) wire n1217_o;
  (* KEEP="TRUE" *) wire n1218_o;
  (* KEEP="TRUE" *) wire n1219_o;
  (* KEEP="TRUE" *) wire n1220_o;
  (* KEEP="TRUE" *) wire n1221_o;
  (* KEEP="TRUE" *) wire n1222_o;
  (* KEEP="TRUE" *) wire n1223_o;
  (* KEEP="TRUE" *) wire n1224_o;
  (* KEEP="TRUE" *) wire n1225_o;
  (* KEEP="TRUE" *) wire n1226_o;
  (* KEEP="TRUE" *) wire n1227_o;
  (* KEEP="TRUE" *) wire n1228_o;
  (* KEEP="TRUE" *) wire n1229_o;
  (* KEEP="TRUE" *) wire n1230_o;
  (* KEEP="TRUE" *) wire n1231_o;
  (* KEEP="TRUE" *) wire n1232_o;
  (* KEEP="TRUE" *) wire n1233_o;
  (* KEEP="TRUE" *) wire n1234_o;
  (* KEEP="TRUE" *) wire n1235_o;
  (* KEEP="TRUE" *) wire n1236_o;
  (* KEEP="TRUE" *) wire n1237_o;
  (* KEEP="TRUE" *) wire n1238_o;
  (* KEEP="TRUE" *) wire n1239_o;
  (* KEEP="TRUE" *) wire n1240_o;
  (* KEEP="TRUE" *) wire n1241_o;
  (* KEEP="TRUE" *) wire n1242_o;
  (* KEEP="TRUE" *) wire n1243_o;
  (* KEEP="TRUE" *) wire n1244_o;
  (* KEEP="TRUE" *) wire n1245_o;
  (* KEEP="TRUE" *) wire n1246_o;
  (* KEEP="TRUE" *) wire n1247_o;
  (* KEEP="TRUE" *) wire n1248_o;
  (* KEEP="TRUE" *) wire n1249_o;
  (* KEEP="TRUE" *) wire n1250_o;
  (* KEEP="TRUE" *) wire n1251_o;
  (* KEEP="TRUE" *) wire n1252_o;
  (* KEEP="TRUE" *) wire n1253_o;
  (* KEEP="TRUE" *) wire n1254_o;
  (* KEEP="TRUE" *) wire n1255_o;
  (* KEEP="TRUE" *) wire n1256_o;
  (* KEEP="TRUE" *) wire n1257_o;
  (* KEEP="TRUE" *) wire n1258_o;
  (* KEEP="TRUE" *) wire n1259_o;
  (* KEEP="TRUE" *) wire n1260_o;
  (* KEEP="TRUE" *) wire n1261_o;
  (* KEEP="TRUE" *) wire n1262_o;
  (* KEEP="TRUE" *) wire n1263_o;
  (* KEEP="TRUE" *) wire n1264_o;
  (* KEEP="TRUE" *) wire n1265_o;
  (* KEEP="TRUE" *) wire n1266_o;
  (* KEEP="TRUE" *) wire n1267_o;
  (* KEEP="TRUE" *) wire n1268_o;
  (* KEEP="TRUE" *) wire n1269_o;
  (* KEEP="TRUE" *) wire n1270_o;
  (* KEEP="TRUE" *) wire n1271_o;
  (* KEEP="TRUE" *) wire n1272_o;
  (* KEEP="TRUE" *) wire n1273_o;
  (* KEEP="TRUE" *) wire n1274_o;
  (* KEEP="TRUE" *) wire n1275_o;
  (* KEEP="TRUE" *) wire n1276_o;
  (* KEEP="TRUE" *) wire n1277_o;
  (* KEEP="TRUE" *) wire n1278_o;
  (* KEEP="TRUE" *) wire n1279_o;
  (* KEEP="TRUE" *) wire n1280_o;
  (* KEEP="TRUE" *) wire n1281_o;
  (* KEEP="TRUE" *) wire n1282_o;
  (* KEEP="TRUE" *) wire n1283_o;
  (* KEEP="TRUE" *) wire n1284_o;
  (* KEEP="TRUE" *) wire n1285_o;
  (* KEEP="TRUE" *) wire n1286_o;
  (* KEEP="TRUE" *) wire n1287_o;
  (* KEEP="TRUE" *) wire n1288_o;
  (* KEEP="TRUE" *) wire n1289_o;
  (* KEEP="TRUE" *) wire n1290_o;
  (* KEEP="TRUE" *) wire n1291_o;
  (* KEEP="TRUE" *) wire n1292_o;
  (* KEEP="TRUE" *) wire n1293_o;
  (* KEEP="TRUE" *) wire n1294_o;
  (* KEEP="TRUE" *) wire n1295_o;
  (* KEEP="TRUE" *) wire n1296_o;
  (* KEEP="TRUE" *) wire n1297_o;
  (* KEEP="TRUE" *) wire n1298_o;
  (* KEEP="TRUE" *) wire n1299_o;
  (* KEEP="TRUE" *) wire n1300_o;
  (* KEEP="TRUE" *) wire n1301_o;
  (* KEEP="TRUE" *) wire n1302_o;
  (* KEEP="TRUE" *) wire n1303_o;
  (* KEEP="TRUE" *) wire n1304_o;
  (* KEEP="TRUE" *) wire n1305_o;
  (* KEEP="TRUE" *) wire n1306_o;
  (* KEEP="TRUE" *) wire n1307_o;
  (* KEEP="TRUE" *) wire n1308_o;
  (* KEEP="TRUE" *) wire n1309_o;
  (* KEEP="TRUE" *) wire n1310_o;
  (* KEEP="TRUE" *) wire n1311_o;
  (* KEEP="TRUE" *) wire n1312_o;
  (* KEEP="TRUE" *) wire n1313_o;
  (* KEEP="TRUE" *) wire n1314_o;
  (* KEEP="TRUE" *) wire n1315_o;
  (* KEEP="TRUE" *) wire n1316_o;
  (* KEEP="TRUE" *) wire n1317_o;
  (* KEEP="TRUE" *) wire n1318_o;
  (* KEEP="TRUE" *) wire n1319_o;
  (* KEEP="TRUE" *) wire n1320_o;
  (* KEEP="TRUE" *) wire n1321_o;
  (* KEEP="TRUE" *) wire n1322_o;
  (* KEEP="TRUE" *) wire n1323_o;
  (* KEEP="TRUE" *) wire n1324_o;
  (* KEEP="TRUE" *) wire n1325_o;
  (* KEEP="TRUE" *) wire n1326_o;
  (* KEEP="TRUE" *) wire n1327_o;
  (* KEEP="TRUE" *) wire n1328_o;
  (* KEEP="TRUE" *) wire n1329_o;
  (* KEEP="TRUE" *) wire n1330_o;
  (* KEEP="TRUE" *) wire n1331_o;
  (* KEEP="TRUE" *) wire n1332_o;
  (* KEEP="TRUE" *) wire n1333_o;
  (* KEEP="TRUE" *) wire n1334_o;
  (* KEEP="TRUE" *) wire n1335_o;
  (* KEEP="TRUE" *) wire n1336_o;
  (* KEEP="TRUE" *) wire n1337_o;
  (* KEEP="TRUE" *) wire n1338_o;
  (* KEEP="TRUE" *) wire n1339_o;
  (* KEEP="TRUE" *) wire n1340_o;
  (* KEEP="TRUE" *) wire n1341_o;
  (* KEEP="TRUE" *) wire n1342_o;
  (* KEEP="TRUE" *) wire n1343_o;
  (* KEEP="TRUE" *) wire n1344_o;
  (* KEEP="TRUE" *) wire n1345_o;
  (* KEEP="TRUE" *) wire n1346_o;
  (* KEEP="TRUE" *) wire n1347_o;
  (* KEEP="TRUE" *) wire n1348_o;
  (* KEEP="TRUE" *) wire n1349_o;
  (* KEEP="TRUE" *) wire n1350_o;
  (* KEEP="TRUE" *) wire n1351_o;
  (* KEEP="TRUE" *) wire n1352_o;
  (* KEEP="TRUE" *) wire n1353_o;
  (* KEEP="TRUE" *) wire n1354_o;
  (* KEEP="TRUE" *) wire n1355_o;
  (* KEEP="TRUE" *) wire n1356_o;
  (* KEEP="TRUE" *) wire n1357_o;
  (* KEEP="TRUE" *) wire n1358_o;
  (* KEEP="TRUE" *) wire n1359_o;
  (* KEEP="TRUE" *) wire n1360_o;
  (* KEEP="TRUE" *) wire n1361_o;
  (* KEEP="TRUE" *) wire n1362_o;
  (* KEEP="TRUE" *) wire n1363_o;
  (* KEEP="TRUE" *) wire n1364_o;
  (* KEEP="TRUE" *) wire n1365_o;
  (* KEEP="TRUE" *) wire n1366_o;
  (* KEEP="TRUE" *) wire n1367_o;
  (* KEEP="TRUE" *) wire n1368_o;
  (* KEEP="TRUE" *) wire n1369_o;
  (* KEEP="TRUE" *) wire n1370_o;
  (* KEEP="TRUE" *) wire n1371_o;
  (* KEEP="TRUE" *) wire n1372_o;
  (* KEEP="TRUE" *) wire n1373_o;
  (* KEEP="TRUE" *) wire n1374_o;
  (* KEEP="TRUE" *) wire n1375_o;
  (* KEEP="TRUE" *) wire n1376_o;
  (* KEEP="TRUE" *) wire n1377_o;
  (* KEEP="TRUE" *) wire n1378_o;
  (* KEEP="TRUE" *) wire n1379_o;
  (* KEEP="TRUE" *) wire n1380_o;
  (* KEEP="TRUE" *) wire n1381_o;
  (* KEEP="TRUE" *) wire n1382_o;
  (* KEEP="TRUE" *) wire n1383_o;
  (* KEEP="TRUE" *) wire n1384_o;
  (* KEEP="TRUE" *) wire n1385_o;
  (* KEEP="TRUE" *) wire n1386_o;
  (* KEEP="TRUE" *) wire n1387_o;
  (* KEEP="TRUE" *) wire n1388_o;
  (* KEEP="TRUE" *) wire n1389_o;
  (* KEEP="TRUE" *) wire n1390_o;
  (* KEEP="TRUE" *) wire n1391_o;
  (* KEEP="TRUE" *) wire n1392_o;
  (* KEEP="TRUE" *) wire n1393_o;
  (* KEEP="TRUE" *) wire n1394_o;
  (* KEEP="TRUE" *) wire n1395_o;
  (* KEEP="TRUE" *) wire n1396_o;
  (* KEEP="TRUE" *) wire n1397_o;
  (* KEEP="TRUE" *) wire n1398_o;
  (* KEEP="TRUE" *) wire n1399_o;
  (* KEEP="TRUE" *) wire n1400_o;
  (* KEEP="TRUE" *) wire n1401_o;
  (* KEEP="TRUE" *) wire n1402_o;
  (* KEEP="TRUE" *) wire n1403_o;
  (* KEEP="TRUE" *) wire n1404_o;
  (* KEEP="TRUE" *) wire n1405_o;
  (* KEEP="TRUE" *) wire n1406_o;
  (* KEEP="TRUE" *) wire n1407_o;
  (* KEEP="TRUE" *) wire n1408_o;
  (* KEEP="TRUE" *) wire n1409_o;
  (* KEEP="TRUE" *) wire n1410_o;
  (* KEEP="TRUE" *) wire n1411_o;
  (* KEEP="TRUE" *) wire n1412_o;
  (* KEEP="TRUE" *) wire n1413_o;
  (* KEEP="TRUE" *) wire n1414_o;
  (* KEEP="TRUE" *) wire n1415_o;
  (* KEEP="TRUE" *) wire n1416_o;
  (* KEEP="TRUE" *) wire n1417_o;
  (* KEEP="TRUE" *) wire n1418_o;
  (* KEEP="TRUE" *) wire n1419_o;
  (* KEEP="TRUE" *) wire n1420_o;
  (* KEEP="TRUE" *) wire n1421_o;
  (* KEEP="TRUE" *) wire n1422_o;
  (* KEEP="TRUE" *) wire n1423_o;
  (* KEEP="TRUE" *) wire n1424_o;
  (* KEEP="TRUE" *) wire n1425_o;
  (* KEEP="TRUE" *) wire n1426_o;
  (* KEEP="TRUE" *) wire n1427_o;
  (* KEEP="TRUE" *) wire n1428_o;
  (* KEEP="TRUE" *) wire n1429_o;
  (* KEEP="TRUE" *) wire n1430_o;
  (* KEEP="TRUE" *) wire n1431_o;
  (* KEEP="TRUE" *) wire n1432_o;
  (* KEEP="TRUE" *) wire n1433_o;
  (* KEEP="TRUE" *) wire n1434_o;
  (* KEEP="TRUE" *) wire n1435_o;
  (* KEEP="TRUE" *) wire n1436_o;
  (* KEEP="TRUE" *) wire n1437_o;
  (* KEEP="TRUE" *) wire n1438_o;
  (* KEEP="TRUE" *) wire n1439_o;
  (* KEEP="TRUE" *) wire n1440_o;
  (* KEEP="TRUE" *) wire n1441_o;
  (* KEEP="TRUE" *) wire n1442_o;
  (* KEEP="TRUE" *) wire n1443_o;
  (* KEEP="TRUE" *) wire n1444_o;
  (* KEEP="TRUE" *) wire n1445_o;
  (* KEEP="TRUE" *) wire n1446_o;
  (* KEEP="TRUE" *) wire n1447_o;
  (* KEEP="TRUE" *) wire n1448_o;
  (* KEEP="TRUE" *) wire n1449_o;
  (* KEEP="TRUE" *) wire n1450_o;
  (* KEEP="TRUE" *) wire n1451_o;
  (* KEEP="TRUE" *) wire n1452_o;
  (* KEEP="TRUE" *) wire n1453_o;
  (* KEEP="TRUE" *) wire n1454_o;
  (* KEEP="TRUE" *) wire n1455_o;
  (* KEEP="TRUE" *) wire n1456_o;
  (* KEEP="TRUE" *) wire n1457_o;
  (* KEEP="TRUE" *) wire n1458_o;
  (* KEEP="TRUE" *) wire n1459_o;
  (* KEEP="TRUE" *) wire n1460_o;
  (* KEEP="TRUE" *) wire n1461_o;
  (* KEEP="TRUE" *) wire n1462_o;
  (* KEEP="TRUE" *) wire n1463_o;
  (* KEEP="TRUE" *) wire n1464_o;
  (* KEEP="TRUE" *) wire n1465_o;
  (* KEEP="TRUE" *) wire n1466_o;
  (* KEEP="TRUE" *) wire n1467_o;
  (* KEEP="TRUE" *) wire n1468_o;
  (* KEEP="TRUE" *) wire n1469_o;
  (* KEEP="TRUE" *) wire n1470_o;
  (* KEEP="TRUE" *) wire n1471_o;
  (* KEEP="TRUE" *) wire n1472_o;
  (* KEEP="TRUE" *) wire n1473_o;
  (* KEEP="TRUE" *) wire n1474_o;
  (* KEEP="TRUE" *) wire n1475_o;
  (* KEEP="TRUE" *) wire n1476_o;
  (* KEEP="TRUE" *) wire n1477_o;
  (* KEEP="TRUE" *) wire n1478_o;
  (* KEEP="TRUE" *) wire n1479_o;
  (* KEEP="TRUE" *) wire n1480_o;
  (* KEEP="TRUE" *) wire n1481_o;
  (* KEEP="TRUE" *) wire n1482_o;
  (* KEEP="TRUE" *) wire n1483_o;
  (* KEEP="TRUE" *) wire n1484_o;
  (* KEEP="TRUE" *) wire n1485_o;
  (* KEEP="TRUE" *) wire n1486_o;
  (* KEEP="TRUE" *) wire n1487_o;
  (* KEEP="TRUE" *) wire n1488_o;
  (* KEEP="TRUE" *) wire n1489_o;
  (* KEEP="TRUE" *) wire n1490_o;
  (* KEEP="TRUE" *) wire n1491_o;
  (* KEEP="TRUE" *) wire n1492_o;
  (* KEEP="TRUE" *) wire n1493_o;
  (* KEEP="TRUE" *) wire n1494_o;
  (* KEEP="TRUE" *) wire n1495_o;
  (* KEEP="TRUE" *) wire n1496_o;
  (* KEEP="TRUE" *) wire n1497_o;
  (* KEEP="TRUE" *) wire n1498_o;
  (* KEEP="TRUE" *) wire n1499_o;
  (* KEEP="TRUE" *) wire n1500_o;
  (* KEEP="TRUE" *) wire n1501_o;
  (* KEEP="TRUE" *) wire n1502_o;
  (* KEEP="TRUE" *) wire n1503_o;
  (* KEEP="TRUE" *) wire n1504_o;
  (* KEEP="TRUE" *) wire n1505_o;
  (* KEEP="TRUE" *) wire n1506_o;
  (* KEEP="TRUE" *) wire n1507_o;
  (* KEEP="TRUE" *) wire n1508_o;
  (* KEEP="TRUE" *) wire n1509_o;
  (* KEEP="TRUE" *) wire n1510_o;
  (* KEEP="TRUE" *) wire n1511_o;
  (* KEEP="TRUE" *) wire n1512_o;
  (* KEEP="TRUE" *) wire n1513_o;
  (* KEEP="TRUE" *) wire n1514_o;
  (* KEEP="TRUE" *) wire n1515_o;
  (* KEEP="TRUE" *) wire n1516_o;
  (* KEEP="TRUE" *) wire n1517_o;
  (* KEEP="TRUE" *) wire n1518_o;
  (* KEEP="TRUE" *) wire n1519_o;
  (* KEEP="TRUE" *) wire n1520_o;
  (* KEEP="TRUE" *) wire n1521_o;
  (* KEEP="TRUE" *) wire n1522_o;
  (* KEEP="TRUE" *) wire n1523_o;
  (* KEEP="TRUE" *) wire n1524_o;
  (* KEEP="TRUE" *) wire n1525_o;
  (* KEEP="TRUE" *) wire n1526_o;
  (* KEEP="TRUE" *) wire n1527_o;
  (* KEEP="TRUE" *) wire n1528_o;
  (* KEEP="TRUE" *) wire n1529_o;
  (* KEEP="TRUE" *) wire n1530_o;
  (* KEEP="TRUE" *) wire n1531_o;
  (* KEEP="TRUE" *) wire n1532_o;
  (* KEEP="TRUE" *) wire [255:0] n1533_o;
  (* KEEP="TRUE" *) wire n1534_o;
  (* KEEP="TRUE" *) wire n1535_o;
  (* KEEP="TRUE" *) wire n1536_o;
  (* KEEP="TRUE" *) wire n1537_o;
  (* KEEP="TRUE" *) wire n1538_o;
  (* KEEP="TRUE" *) wire n1539_o;
  (* KEEP="TRUE" *) wire n1540_o;
  (* KEEP="TRUE" *) wire n1541_o;
  (* KEEP="TRUE" *) wire n1542_o;
  (* KEEP="TRUE" *) wire n1543_o;
  (* KEEP="TRUE" *) wire n1544_o;
  (* KEEP="TRUE" *) wire n1545_o;
  (* KEEP="TRUE" *) wire n1546_o;
  (* KEEP="TRUE" *) wire n1547_o;
  (* KEEP="TRUE" *) wire n1548_o;
  (* KEEP="TRUE" *) wire n1549_o;
  (* KEEP="TRUE" *) wire n1550_o;
  (* KEEP="TRUE" *) wire n1551_o;
  (* KEEP="TRUE" *) wire n1552_o;
  (* KEEP="TRUE" *) wire n1553_o;
  (* KEEP="TRUE" *) wire n1554_o;
  (* KEEP="TRUE" *) wire n1555_o;
  (* KEEP="TRUE" *) wire n1556_o;
  (* KEEP="TRUE" *) wire n1557_o;
  (* KEEP="TRUE" *) wire n1558_o;
  (* KEEP="TRUE" *) wire n1559_o;
  (* KEEP="TRUE" *) wire n1560_o;
  (* KEEP="TRUE" *) wire n1561_o;
  (* KEEP="TRUE" *) wire n1562_o;
  (* KEEP="TRUE" *) wire n1563_o;
  (* KEEP="TRUE" *) wire n1564_o;
  (* KEEP="TRUE" *) wire n1565_o;
  (* KEEP="TRUE" *) wire n1566_o;
  (* KEEP="TRUE" *) wire n1567_o;
  (* KEEP="TRUE" *) wire n1568_o;
  (* KEEP="TRUE" *) wire n1569_o;
  (* KEEP="TRUE" *) wire n1570_o;
  (* KEEP="TRUE" *) wire n1571_o;
  (* KEEP="TRUE" *) wire n1572_o;
  (* KEEP="TRUE" *) wire n1573_o;
  (* KEEP="TRUE" *) wire n1574_o;
  (* KEEP="TRUE" *) wire n1575_o;
  (* KEEP="TRUE" *) wire n1576_o;
  (* KEEP="TRUE" *) wire n1577_o;
  (* KEEP="TRUE" *) wire n1578_o;
  (* KEEP="TRUE" *) wire n1579_o;
  (* KEEP="TRUE" *) wire n1580_o;
  (* KEEP="TRUE" *) wire n1581_o;
  (* KEEP="TRUE" *) wire n1582_o;
  (* KEEP="TRUE" *) wire n1583_o;
  (* KEEP="TRUE" *) wire n1584_o;
  (* KEEP="TRUE" *) wire n1585_o;
  (* KEEP="TRUE" *) wire n1586_o;
  (* KEEP="TRUE" *) wire n1587_o;
  (* KEEP="TRUE" *) wire n1588_o;
  (* KEEP="TRUE" *) wire n1589_o;
  (* KEEP="TRUE" *) wire n1590_o;
  (* KEEP="TRUE" *) wire n1591_o;
  (* KEEP="TRUE" *) wire n1592_o;
  (* KEEP="TRUE" *) wire n1593_o;
  (* KEEP="TRUE" *) wire n1594_o;
  (* KEEP="TRUE" *) wire n1595_o;
  (* KEEP="TRUE" *) wire n1596_o;
  (* KEEP="TRUE" *) wire n1597_o;
  (* KEEP="TRUE" *) wire n1598_o;
  (* KEEP="TRUE" *) wire n1599_o;
  (* KEEP="TRUE" *) wire n1600_o;
  (* KEEP="TRUE" *) wire n1601_o;
  (* KEEP="TRUE" *) wire n1602_o;
  (* KEEP="TRUE" *) wire n1603_o;
  (* KEEP="TRUE" *) wire n1604_o;
  (* KEEP="TRUE" *) wire n1605_o;
  (* KEEP="TRUE" *) wire n1606_o;
  (* KEEP="TRUE" *) wire n1607_o;
  (* KEEP="TRUE" *) wire n1608_o;
  (* KEEP="TRUE" *) wire n1609_o;
  (* KEEP="TRUE" *) wire n1610_o;
  (* KEEP="TRUE" *) wire n1611_o;
  (* KEEP="TRUE" *) wire n1612_o;
  (* KEEP="TRUE" *) wire n1613_o;
  (* KEEP="TRUE" *) wire n1614_o;
  (* KEEP="TRUE" *) wire n1615_o;
  (* KEEP="TRUE" *) wire n1616_o;
  (* KEEP="TRUE" *) wire n1617_o;
  (* KEEP="TRUE" *) wire n1618_o;
  (* KEEP="TRUE" *) wire n1619_o;
  (* KEEP="TRUE" *) wire n1620_o;
  (* KEEP="TRUE" *) wire n1621_o;
  (* KEEP="TRUE" *) wire n1622_o;
  (* KEEP="TRUE" *) wire n1623_o;
  (* KEEP="TRUE" *) wire n1624_o;
  (* KEEP="TRUE" *) wire n1625_o;
  (* KEEP="TRUE" *) wire n1626_o;
  (* KEEP="TRUE" *) wire n1627_o;
  (* KEEP="TRUE" *) wire n1628_o;
  (* KEEP="TRUE" *) wire n1629_o;
  (* KEEP="TRUE" *) wire n1630_o;
  (* KEEP="TRUE" *) wire n1631_o;
  (* KEEP="TRUE" *) wire n1632_o;
  (* KEEP="TRUE" *) wire n1633_o;
  (* KEEP="TRUE" *) wire n1634_o;
  (* KEEP="TRUE" *) wire n1635_o;
  (* KEEP="TRUE" *) wire n1636_o;
  (* KEEP="TRUE" *) wire n1637_o;
  (* KEEP="TRUE" *) wire n1638_o;
  (* KEEP="TRUE" *) wire n1639_o;
  (* KEEP="TRUE" *) wire n1640_o;
  (* KEEP="TRUE" *) wire n1641_o;
  (* KEEP="TRUE" *) wire n1642_o;
  (* KEEP="TRUE" *) wire n1643_o;
  (* KEEP="TRUE" *) wire n1644_o;
  (* KEEP="TRUE" *) wire n1645_o;
  (* KEEP="TRUE" *) wire n1646_o;
  (* KEEP="TRUE" *) wire n1647_o;
  (* KEEP="TRUE" *) wire n1648_o;
  (* KEEP="TRUE" *) wire n1649_o;
  (* KEEP="TRUE" *) wire n1650_o;
  (* KEEP="TRUE" *) wire n1651_o;
  (* KEEP="TRUE" *) wire n1652_o;
  (* KEEP="TRUE" *) wire n1653_o;
  (* KEEP="TRUE" *) wire n1654_o;
  (* KEEP="TRUE" *) wire n1655_o;
  (* KEEP="TRUE" *) wire n1656_o;
  (* KEEP="TRUE" *) wire n1657_o;
  (* KEEP="TRUE" *) wire n1658_o;
  (* KEEP="TRUE" *) wire n1659_o;
  (* KEEP="TRUE" *) wire n1660_o;
  (* KEEP="TRUE" *) wire n1661_o;
  (* KEEP="TRUE" *) wire n1662_o;
  (* KEEP="TRUE" *) wire n1663_o;
  (* KEEP="TRUE" *) wire n1664_o;
  (* KEEP="TRUE" *) wire n1665_o;
  (* KEEP="TRUE" *) wire n1666_o;
  (* KEEP="TRUE" *) wire n1667_o;
  (* KEEP="TRUE" *) wire n1668_o;
  (* KEEP="TRUE" *) wire n1669_o;
  (* KEEP="TRUE" *) wire n1670_o;
  (* KEEP="TRUE" *) wire n1671_o;
  (* KEEP="TRUE" *) wire n1672_o;
  (* KEEP="TRUE" *) wire n1673_o;
  (* KEEP="TRUE" *) wire n1674_o;
  (* KEEP="TRUE" *) wire n1675_o;
  (* KEEP="TRUE" *) wire n1676_o;
  (* KEEP="TRUE" *) wire n1677_o;
  (* KEEP="TRUE" *) wire n1678_o;
  (* KEEP="TRUE" *) wire n1679_o;
  (* KEEP="TRUE" *) wire n1680_o;
  (* KEEP="TRUE" *) wire n1681_o;
  (* KEEP="TRUE" *) wire n1682_o;
  (* KEEP="TRUE" *) wire n1683_o;
  (* KEEP="TRUE" *) wire n1684_o;
  (* KEEP="TRUE" *) wire n1685_o;
  (* KEEP="TRUE" *) wire n1686_o;
  (* KEEP="TRUE" *) wire n1687_o;
  (* KEEP="TRUE" *) wire n1688_o;
  (* KEEP="TRUE" *) wire n1689_o;
  (* KEEP="TRUE" *) wire n1690_o;
  (* KEEP="TRUE" *) wire n1691_o;
  (* KEEP="TRUE" *) wire n1692_o;
  (* KEEP="TRUE" *) wire n1693_o;
  (* KEEP="TRUE" *) wire n1694_o;
  (* KEEP="TRUE" *) wire n1695_o;
  (* KEEP="TRUE" *) wire n1696_o;
  (* KEEP="TRUE" *) wire n1697_o;
  (* KEEP="TRUE" *) wire n1698_o;
  (* KEEP="TRUE" *) wire n1699_o;
  (* KEEP="TRUE" *) wire n1700_o;
  (* KEEP="TRUE" *) wire n1701_o;
  (* KEEP="TRUE" *) wire n1702_o;
  (* KEEP="TRUE" *) wire n1703_o;
  (* KEEP="TRUE" *) wire n1704_o;
  (* KEEP="TRUE" *) wire n1705_o;
  (* KEEP="TRUE" *) wire n1706_o;
  (* KEEP="TRUE" *) wire n1707_o;
  (* KEEP="TRUE" *) wire n1708_o;
  (* KEEP="TRUE" *) wire n1709_o;
  (* KEEP="TRUE" *) wire n1710_o;
  (* KEEP="TRUE" *) wire n1711_o;
  (* KEEP="TRUE" *) wire n1712_o;
  (* KEEP="TRUE" *) wire n1713_o;
  (* KEEP="TRUE" *) wire n1714_o;
  (* KEEP="TRUE" *) wire n1715_o;
  (* KEEP="TRUE" *) wire n1716_o;
  (* KEEP="TRUE" *) wire n1717_o;
  (* KEEP="TRUE" *) wire n1718_o;
  (* KEEP="TRUE" *) wire n1719_o;
  (* KEEP="TRUE" *) wire n1720_o;
  (* KEEP="TRUE" *) wire n1721_o;
  (* KEEP="TRUE" *) wire n1722_o;
  (* KEEP="TRUE" *) wire n1723_o;
  (* KEEP="TRUE" *) wire n1724_o;
  (* KEEP="TRUE" *) wire n1725_o;
  (* KEEP="TRUE" *) wire n1726_o;
  (* KEEP="TRUE" *) wire n1727_o;
  (* KEEP="TRUE" *) wire n1728_o;
  (* KEEP="TRUE" *) wire n1729_o;
  (* KEEP="TRUE" *) wire n1730_o;
  (* KEEP="TRUE" *) wire n1731_o;
  (* KEEP="TRUE" *) wire n1732_o;
  (* KEEP="TRUE" *) wire n1733_o;
  (* KEEP="TRUE" *) wire n1734_o;
  (* KEEP="TRUE" *) wire n1735_o;
  (* KEEP="TRUE" *) wire n1736_o;
  (* KEEP="TRUE" *) wire n1737_o;
  (* KEEP="TRUE" *) wire n1738_o;
  (* KEEP="TRUE" *) wire n1739_o;
  (* KEEP="TRUE" *) wire n1740_o;
  (* KEEP="TRUE" *) wire n1741_o;
  (* KEEP="TRUE" *) wire n1742_o;
  (* KEEP="TRUE" *) wire n1743_o;
  (* KEEP="TRUE" *) wire n1744_o;
  (* KEEP="TRUE" *) wire n1745_o;
  (* KEEP="TRUE" *) wire n1746_o;
  (* KEEP="TRUE" *) wire n1747_o;
  (* KEEP="TRUE" *) wire n1748_o;
  (* KEEP="TRUE" *) wire n1749_o;
  (* KEEP="TRUE" *) wire n1750_o;
  (* KEEP="TRUE" *) wire n1751_o;
  (* KEEP="TRUE" *) wire n1752_o;
  (* KEEP="TRUE" *) wire n1753_o;
  (* KEEP="TRUE" *) wire n1754_o;
  (* KEEP="TRUE" *) wire n1755_o;
  (* KEEP="TRUE" *) wire n1756_o;
  (* KEEP="TRUE" *) wire n1757_o;
  (* KEEP="TRUE" *) wire n1758_o;
  (* KEEP="TRUE" *) wire n1759_o;
  (* KEEP="TRUE" *) wire n1760_o;
  (* KEEP="TRUE" *) wire n1761_o;
  (* KEEP="TRUE" *) wire n1762_o;
  (* KEEP="TRUE" *) wire n1763_o;
  (* KEEP="TRUE" *) wire n1764_o;
  (* KEEP="TRUE" *) wire n1765_o;
  (* KEEP="TRUE" *) wire n1766_o;
  (* KEEP="TRUE" *) wire n1767_o;
  (* KEEP="TRUE" *) wire n1768_o;
  (* KEEP="TRUE" *) wire n1769_o;
  (* KEEP="TRUE" *) wire n1770_o;
  (* KEEP="TRUE" *) wire n1771_o;
  (* KEEP="TRUE" *) wire n1772_o;
  (* KEEP="TRUE" *) wire n1773_o;
  (* KEEP="TRUE" *) wire n1774_o;
  (* KEEP="TRUE" *) wire n1775_o;
  (* KEEP="TRUE" *) wire n1776_o;
  (* KEEP="TRUE" *) wire n1777_o;
  (* KEEP="TRUE" *) wire n1778_o;
  (* KEEP="TRUE" *) wire n1779_o;
  (* KEEP="TRUE" *) wire n1780_o;
  (* KEEP="TRUE" *) wire n1781_o;
  (* KEEP="TRUE" *) wire n1782_o;
  (* KEEP="TRUE" *) wire n1783_o;
  (* KEEP="TRUE" *) wire n1784_o;
  (* KEEP="TRUE" *) wire n1785_o;
  (* KEEP="TRUE" *) wire n1786_o;
  (* KEEP="TRUE" *) wire n1787_o;
  (* KEEP="TRUE" *) wire n1788_o;
  (* KEEP="TRUE" *) wire n1789_o;
  (* KEEP="TRUE" *) wire n1790_o;
  (* KEEP="TRUE" *) wire n1791_o;
  (* KEEP="TRUE" *) wire n1792_o;
  (* KEEP="TRUE" *) wire n1793_o;
  (* KEEP="TRUE" *) wire n1794_o;
  (* KEEP="TRUE" *) wire n1795_o;
  (* KEEP="TRUE" *) wire n1796_o;
  (* KEEP="TRUE" *) wire n1797_o;
  (* KEEP="TRUE" *) wire n1798_o;
  (* KEEP="TRUE" *) wire n1799_o;
  (* KEEP="TRUE" *) wire n1800_o;
  (* KEEP="TRUE" *) wire n1801_o;
  (* KEEP="TRUE" *) wire n1802_o;
  (* KEEP="TRUE" *) wire n1803_o;
  (* KEEP="TRUE" *) wire n1804_o;
  (* KEEP="TRUE" *) wire n1805_o;
  (* KEEP="TRUE" *) wire n1806_o;
  (* KEEP="TRUE" *) wire n1807_o;
  (* KEEP="TRUE" *) wire n1808_o;
  (* KEEP="TRUE" *) wire n1809_o;
  (* KEEP="TRUE" *) wire n1810_o;
  (* KEEP="TRUE" *) wire n1811_o;
  (* KEEP="TRUE" *) wire n1812_o;
  (* KEEP="TRUE" *) wire n1813_o;
  (* KEEP="TRUE" *) wire n1814_o;
  (* KEEP="TRUE" *) wire n1815_o;
  (* KEEP="TRUE" *) wire n1816_o;
  (* KEEP="TRUE" *) wire n1817_o;
  (* KEEP="TRUE" *) wire n1818_o;
  (* KEEP="TRUE" *) wire n1819_o;
  (* KEEP="TRUE" *) wire n1820_o;
  (* KEEP="TRUE" *) wire n1821_o;
  (* KEEP="TRUE" *) wire n1822_o;
  (* KEEP="TRUE" *) wire n1823_o;
  (* KEEP="TRUE" *) wire n1824_o;
  (* KEEP="TRUE" *) wire n1825_o;
  (* KEEP="TRUE" *) wire n1826_o;
  (* KEEP="TRUE" *) wire n1827_o;
  (* KEEP="TRUE" *) wire n1828_o;
  (* KEEP="TRUE" *) wire n1829_o;
  (* KEEP="TRUE" *) wire n1830_o;
  (* KEEP="TRUE" *) wire n1831_o;
  (* KEEP="TRUE" *) wire n1832_o;
  (* KEEP="TRUE" *) wire n1833_o;
  (* KEEP="TRUE" *) wire n1834_o;
  (* KEEP="TRUE" *) wire n1835_o;
  (* KEEP="TRUE" *) wire n1836_o;
  (* KEEP="TRUE" *) wire n1837_o;
  (* KEEP="TRUE" *) wire n1838_o;
  (* KEEP="TRUE" *) wire n1839_o;
  (* KEEP="TRUE" *) wire n1840_o;
  (* KEEP="TRUE" *) wire n1841_o;
  (* KEEP="TRUE" *) wire n1842_o;
  (* KEEP="TRUE" *) wire n1843_o;
  (* KEEP="TRUE" *) wire n1844_o;
  (* KEEP="TRUE" *) wire n1845_o;
  (* KEEP="TRUE" *) wire n1846_o;
  (* KEEP="TRUE" *) wire n1847_o;
  (* KEEP="TRUE" *) wire n1848_o;
  (* KEEP="TRUE" *) wire n1849_o;
  (* KEEP="TRUE" *) wire n1850_o;
  (* KEEP="TRUE" *) wire n1851_o;
  (* KEEP="TRUE" *) wire n1852_o;
  (* KEEP="TRUE" *) wire n1853_o;
  (* KEEP="TRUE" *) wire n1854_o;
  (* KEEP="TRUE" *) wire n1855_o;
  (* KEEP="TRUE" *) wire n1856_o;
  (* KEEP="TRUE" *) wire n1857_o;
  (* KEEP="TRUE" *) wire n1858_o;
  (* KEEP="TRUE" *) wire n1859_o;
  (* KEEP="TRUE" *) wire n1860_o;
  (* KEEP="TRUE" *) wire n1861_o;
  (* KEEP="TRUE" *) wire n1862_o;
  (* KEEP="TRUE" *) wire n1863_o;
  (* KEEP="TRUE" *) wire n1864_o;
  (* KEEP="TRUE" *) wire n1865_o;
  (* KEEP="TRUE" *) wire n1866_o;
  (* KEEP="TRUE" *) wire n1867_o;
  (* KEEP="TRUE" *) wire n1868_o;
  (* KEEP="TRUE" *) wire n1869_o;
  (* KEEP="TRUE" *) wire n1870_o;
  (* KEEP="TRUE" *) wire n1871_o;
  (* KEEP="TRUE" *) wire n1872_o;
  (* KEEP="TRUE" *) wire n1873_o;
  (* KEEP="TRUE" *) wire n1874_o;
  (* KEEP="TRUE" *) wire n1875_o;
  (* KEEP="TRUE" *) wire n1876_o;
  (* KEEP="TRUE" *) wire n1877_o;
  (* KEEP="TRUE" *) wire n1878_o;
  (* KEEP="TRUE" *) wire n1879_o;
  (* KEEP="TRUE" *) wire n1880_o;
  (* KEEP="TRUE" *) wire n1881_o;
  (* KEEP="TRUE" *) wire n1882_o;
  (* KEEP="TRUE" *) wire n1883_o;
  (* KEEP="TRUE" *) wire n1884_o;
  (* KEEP="TRUE" *) wire n1885_o;
  (* KEEP="TRUE" *) wire n1886_o;
  (* KEEP="TRUE" *) wire n1887_o;
  (* KEEP="TRUE" *) wire n1888_o;
  (* KEEP="TRUE" *) wire n1889_o;
  (* KEEP="TRUE" *) wire n1890_o;
  (* KEEP="TRUE" *) wire n1891_o;
  (* KEEP="TRUE" *) wire n1892_o;
  (* KEEP="TRUE" *) wire n1893_o;
  (* KEEP="TRUE" *) wire n1894_o;
  (* KEEP="TRUE" *) wire n1895_o;
  (* KEEP="TRUE" *) wire n1896_o;
  (* KEEP="TRUE" *) wire n1897_o;
  (* KEEP="TRUE" *) wire n1898_o;
  (* KEEP="TRUE" *) wire n1899_o;
  (* KEEP="TRUE" *) wire n1900_o;
  (* KEEP="TRUE" *) wire n1901_o;
  (* KEEP="TRUE" *) wire n1902_o;
  (* KEEP="TRUE" *) wire n1903_o;
  (* KEEP="TRUE" *) wire n1904_o;
  (* KEEP="TRUE" *) wire n1905_o;
  (* KEEP="TRUE" *) wire n1906_o;
  (* KEEP="TRUE" *) wire n1907_o;
  (* KEEP="TRUE" *) wire n1908_o;
  (* KEEP="TRUE" *) wire n1909_o;
  (* KEEP="TRUE" *) wire n1910_o;
  (* KEEP="TRUE" *) wire n1911_o;
  (* KEEP="TRUE" *) wire n1912_o;
  (* KEEP="TRUE" *) wire n1913_o;
  (* KEEP="TRUE" *) wire n1914_o;
  (* KEEP="TRUE" *) wire n1915_o;
  (* KEEP="TRUE" *) wire n1916_o;
  (* KEEP="TRUE" *) wire n1917_o;
  (* KEEP="TRUE" *) wire n1918_o;
  (* KEEP="TRUE" *) wire n1919_o;
  (* KEEP="TRUE" *) wire n1920_o;
  (* KEEP="TRUE" *) wire n1921_o;
  (* KEEP="TRUE" *) wire n1922_o;
  (* KEEP="TRUE" *) wire n1923_o;
  (* KEEP="TRUE" *) wire n1924_o;
  (* KEEP="TRUE" *) wire n1925_o;
  (* KEEP="TRUE" *) wire n1926_o;
  (* KEEP="TRUE" *) wire n1927_o;
  (* KEEP="TRUE" *) wire n1928_o;
  (* KEEP="TRUE" *) wire n1929_o;
  (* KEEP="TRUE" *) wire n1930_o;
  (* KEEP="TRUE" *) wire n1931_o;
  (* KEEP="TRUE" *) wire n1932_o;
  (* KEEP="TRUE" *) wire n1933_o;
  (* KEEP="TRUE" *) wire n1934_o;
  (* KEEP="TRUE" *) wire n1935_o;
  (* KEEP="TRUE" *) wire n1936_o;
  (* KEEP="TRUE" *) wire n1937_o;
  (* KEEP="TRUE" *) wire n1938_o;
  (* KEEP="TRUE" *) wire n1939_o;
  (* KEEP="TRUE" *) wire n1940_o;
  (* KEEP="TRUE" *) wire n1941_o;
  (* KEEP="TRUE" *) wire n1942_o;
  (* KEEP="TRUE" *) wire n1943_o;
  (* KEEP="TRUE" *) wire n1944_o;
  (* KEEP="TRUE" *) wire n1945_o;
  (* KEEP="TRUE" *) wire n1946_o;
  (* KEEP="TRUE" *) wire n1947_o;
  (* KEEP="TRUE" *) wire n1948_o;
  (* KEEP="TRUE" *) wire n1949_o;
  (* KEEP="TRUE" *) wire n1950_o;
  (* KEEP="TRUE" *) wire n1951_o;
  (* KEEP="TRUE" *) wire n1952_o;
  (* KEEP="TRUE" *) wire n1953_o;
  (* KEEP="TRUE" *) wire n1954_o;
  (* KEEP="TRUE" *) wire n1955_o;
  (* KEEP="TRUE" *) wire n1956_o;
  (* KEEP="TRUE" *) wire n1957_o;
  (* KEEP="TRUE" *) wire n1958_o;
  (* KEEP="TRUE" *) wire n1959_o;
  (* KEEP="TRUE" *) wire n1960_o;
  (* KEEP="TRUE" *) wire n1961_o;
  (* KEEP="TRUE" *) wire n1962_o;
  (* KEEP="TRUE" *) wire n1963_o;
  (* KEEP="TRUE" *) wire n1964_o;
  (* KEEP="TRUE" *) wire n1965_o;
  (* KEEP="TRUE" *) wire n1966_o;
  (* KEEP="TRUE" *) wire n1967_o;
  (* KEEP="TRUE" *) wire n1968_o;
  (* KEEP="TRUE" *) wire n1969_o;
  (* KEEP="TRUE" *) wire n1970_o;
  (* KEEP="TRUE" *) wire n1971_o;
  (* KEEP="TRUE" *) wire n1972_o;
  (* KEEP="TRUE" *) wire n1973_o;
  (* KEEP="TRUE" *) wire n1974_o;
  (* KEEP="TRUE" *) wire n1975_o;
  (* KEEP="TRUE" *) wire n1976_o;
  (* KEEP="TRUE" *) wire n1977_o;
  (* KEEP="TRUE" *) wire n1978_o;
  (* KEEP="TRUE" *) wire n1979_o;
  (* KEEP="TRUE" *) wire n1980_o;
  (* KEEP="TRUE" *) wire n1981_o;
  (* KEEP="TRUE" *) wire n1982_o;
  (* KEEP="TRUE" *) wire n1983_o;
  (* KEEP="TRUE" *) wire n1984_o;
  (* KEEP="TRUE" *) wire n1985_o;
  (* KEEP="TRUE" *) wire n1986_o;
  (* KEEP="TRUE" *) wire n1987_o;
  (* KEEP="TRUE" *) wire n1988_o;
  (* KEEP="TRUE" *) wire n1989_o;
  (* KEEP="TRUE" *) wire n1990_o;
  (* KEEP="TRUE" *) wire n1991_o;
  (* KEEP="TRUE" *) wire n1992_o;
  (* KEEP="TRUE" *) wire n1993_o;
  (* KEEP="TRUE" *) wire n1994_o;
  (* KEEP="TRUE" *) wire n1995_o;
  (* KEEP="TRUE" *) wire n1996_o;
  (* KEEP="TRUE" *) wire n1997_o;
  (* KEEP="TRUE" *) wire n1998_o;
  (* KEEP="TRUE" *) wire n1999_o;
  (* KEEP="TRUE" *) wire n2000_o;
  (* KEEP="TRUE" *) wire n2001_o;
  (* KEEP="TRUE" *) wire n2002_o;
  (* KEEP="TRUE" *) wire n2003_o;
  (* KEEP="TRUE" *) wire n2004_o;
  (* KEEP="TRUE" *) wire n2005_o;
  (* KEEP="TRUE" *) wire n2006_o;
  (* KEEP="TRUE" *) wire n2007_o;
  (* KEEP="TRUE" *) wire n2008_o;
  (* KEEP="TRUE" *) wire n2009_o;
  (* KEEP="TRUE" *) wire n2010_o;
  (* KEEP="TRUE" *) wire n2011_o;
  (* KEEP="TRUE" *) wire n2012_o;
  (* KEEP="TRUE" *) wire n2013_o;
  (* KEEP="TRUE" *) wire n2014_o;
  (* KEEP="TRUE" *) wire n2015_o;
  (* KEEP="TRUE" *) wire n2016_o;
  (* KEEP="TRUE" *) wire n2017_o;
  (* KEEP="TRUE" *) wire n2018_o;
  (* KEEP="TRUE" *) wire n2019_o;
  (* KEEP="TRUE" *) wire n2020_o;
  (* KEEP="TRUE" *) wire n2021_o;
  (* KEEP="TRUE" *) wire n2022_o;
  (* KEEP="TRUE" *) wire n2023_o;
  (* KEEP="TRUE" *) wire n2024_o;
  (* KEEP="TRUE" *) wire n2025_o;
  (* KEEP="TRUE" *) wire n2026_o;
  (* KEEP="TRUE" *) wire n2027_o;
  (* KEEP="TRUE" *) wire n2028_o;
  (* KEEP="TRUE" *) wire n2029_o;
  (* KEEP="TRUE" *) wire n2030_o;
  (* KEEP="TRUE" *) wire n2031_o;
  (* KEEP="TRUE" *) wire n2032_o;
  (* KEEP="TRUE" *) wire n2033_o;
  (* KEEP="TRUE" *) wire n2034_o;
  (* KEEP="TRUE" *) wire n2035_o;
  (* KEEP="TRUE" *) wire n2036_o;
  (* KEEP="TRUE" *) wire n2037_o;
  (* KEEP="TRUE" *) wire n2038_o;
  (* KEEP="TRUE" *) wire n2039_o;
  (* KEEP="TRUE" *) wire n2040_o;
  (* KEEP="TRUE" *) wire n2041_o;
  (* KEEP="TRUE" *) wire n2042_o;
  (* KEEP="TRUE" *) wire n2043_o;
  (* KEEP="TRUE" *) wire n2044_o;
  (* KEEP="TRUE" *) wire n2045_o;
  (* KEEP="TRUE" *) wire n2046_o;
  (* KEEP="TRUE" *) wire n2047_o;
  (* KEEP="TRUE" *) wire n2048_o;
  (* KEEP="TRUE" *) wire n2049_o;
  (* KEEP="TRUE" *) wire n2050_o;
  (* KEEP="TRUE" *) wire n2051_o;
  (* KEEP="TRUE" *) wire n2052_o;
  (* KEEP="TRUE" *) wire n2053_o;
  (* KEEP="TRUE" *) wire n2054_o;
  (* KEEP="TRUE" *) wire n2055_o;
  (* KEEP="TRUE" *) wire n2056_o;
  (* KEEP="TRUE" *) wire n2057_o;
  (* KEEP="TRUE" *) wire n2058_o;
  (* KEEP="TRUE" *) wire n2059_o;
  (* KEEP="TRUE" *) wire n2060_o;
  (* KEEP="TRUE" *) wire n2061_o;
  (* KEEP="TRUE" *) wire n2062_o;
  (* KEEP="TRUE" *) wire n2063_o;
  (* KEEP="TRUE" *) wire n2064_o;
  (* KEEP="TRUE" *) wire n2065_o;
  (* KEEP="TRUE" *) wire n2066_o;
  (* KEEP="TRUE" *) wire n2067_o;
  (* KEEP="TRUE" *) wire n2068_o;
  (* KEEP="TRUE" *) wire n2069_o;
  (* KEEP="TRUE" *) wire n2070_o;
  (* KEEP="TRUE" *) wire n2071_o;
  (* KEEP="TRUE" *) wire n2072_o;
  (* KEEP="TRUE" *) wire n2073_o;
  (* KEEP="TRUE" *) wire n2074_o;
  (* KEEP="TRUE" *) wire n2075_o;
  (* KEEP="TRUE" *) wire n2076_o;
  (* KEEP="TRUE" *) wire n2077_o;
  (* KEEP="TRUE" *) wire n2078_o;
  (* KEEP="TRUE" *) wire n2079_o;
  (* KEEP="TRUE" *) wire n2080_o;
  (* KEEP="TRUE" *) wire n2081_o;
  (* KEEP="TRUE" *) wire n2082_o;
  (* KEEP="TRUE" *) wire n2083_o;
  (* KEEP="TRUE" *) wire n2084_o;
  (* KEEP="TRUE" *) wire n2085_o;
  (* KEEP="TRUE" *) wire n2086_o;
  (* KEEP="TRUE" *) wire n2087_o;
  (* KEEP="TRUE" *) wire n2088_o;
  (* KEEP="TRUE" *) wire n2089_o;
  (* KEEP="TRUE" *) wire n2090_o;
  (* KEEP="TRUE" *) wire n2091_o;
  (* KEEP="TRUE" *) wire n2092_o;
  (* KEEP="TRUE" *) wire n2093_o;
  (* KEEP="TRUE" *) wire n2094_o;
  (* KEEP="TRUE" *) wire n2095_o;
  (* KEEP="TRUE" *) wire n2096_o;
  (* KEEP="TRUE" *) wire n2097_o;
  (* KEEP="TRUE" *) wire n2098_o;
  (* KEEP="TRUE" *) wire n2099_o;
  (* KEEP="TRUE" *) wire n2100_o;
  (* KEEP="TRUE" *) wire n2101_o;
  (* KEEP="TRUE" *) wire n2102_o;
  (* KEEP="TRUE" *) wire n2103_o;
  (* KEEP="TRUE" *) wire n2104_o;
  (* KEEP="TRUE" *) wire n2105_o;
  (* KEEP="TRUE" *) wire n2106_o;
  (* KEEP="TRUE" *) wire n2107_o;
  (* KEEP="TRUE" *) wire n2108_o;
  (* KEEP="TRUE" *) wire n2109_o;
  (* KEEP="TRUE" *) wire n2110_o;
  (* KEEP="TRUE" *) wire n2111_o;
  (* KEEP="TRUE" *) wire n2112_o;
  (* KEEP="TRUE" *) wire n2113_o;
  (* KEEP="TRUE" *) wire n2114_o;
  (* KEEP="TRUE" *) wire n2115_o;
  (* KEEP="TRUE" *) wire n2116_o;
  (* KEEP="TRUE" *) wire n2117_o;
  (* KEEP="TRUE" *) wire n2118_o;
  (* KEEP="TRUE" *) wire n2119_o;
  (* KEEP="TRUE" *) wire n2120_o;
  (* KEEP="TRUE" *) wire n2121_o;
  (* KEEP="TRUE" *) wire n2122_o;
  (* KEEP="TRUE" *) wire n2123_o;
  (* KEEP="TRUE" *) wire n2124_o;
  (* KEEP="TRUE" *) wire n2125_o;
  (* KEEP="TRUE" *) wire n2126_o;
  (* KEEP="TRUE" *) wire n2127_o;
  (* KEEP="TRUE" *) wire n2128_o;
  (* KEEP="TRUE" *) wire n2129_o;
  (* KEEP="TRUE" *) wire n2130_o;
  (* KEEP="TRUE" *) wire n2131_o;
  (* KEEP="TRUE" *) wire n2132_o;
  (* KEEP="TRUE" *) wire n2133_o;
  (* KEEP="TRUE" *) wire n2134_o;
  (* KEEP="TRUE" *) wire n2135_o;
  (* KEEP="TRUE" *) wire n2136_o;
  (* KEEP="TRUE" *) wire n2137_o;
  (* KEEP="TRUE" *) wire n2138_o;
  (* KEEP="TRUE" *) wire n2139_o;
  (* KEEP="TRUE" *) wire n2140_o;
  (* KEEP="TRUE" *) wire n2141_o;
  (* KEEP="TRUE" *) wire n2142_o;
  (* KEEP="TRUE" *) wire n2143_o;
  (* KEEP="TRUE" *) wire n2144_o;
  (* KEEP="TRUE" *) wire n2145_o;
  (* KEEP="TRUE" *) wire n2146_o;
  (* KEEP="TRUE" *) wire n2147_o;
  (* KEEP="TRUE" *) wire n2148_o;
  (* KEEP="TRUE" *) wire n2149_o;
  (* KEEP="TRUE" *) wire n2150_o;
  (* KEEP="TRUE" *) wire n2151_o;
  (* KEEP="TRUE" *) wire n2152_o;
  (* KEEP="TRUE" *) wire n2153_o;
  (* KEEP="TRUE" *) wire n2154_o;
  (* KEEP="TRUE" *) wire n2155_o;
  (* KEEP="TRUE" *) wire n2156_o;
  (* KEEP="TRUE" *) wire n2157_o;
  (* KEEP="TRUE" *) wire n2158_o;
  (* KEEP="TRUE" *) wire n2159_o;
  (* KEEP="TRUE" *) wire n2160_o;
  (* KEEP="TRUE" *) wire n2161_o;
  (* KEEP="TRUE" *) wire n2162_o;
  (* KEEP="TRUE" *) wire n2163_o;
  (* KEEP="TRUE" *) wire n2164_o;
  (* KEEP="TRUE" *) wire n2165_o;
  (* KEEP="TRUE" *) wire n2166_o;
  (* KEEP="TRUE" *) wire n2167_o;
  (* KEEP="TRUE" *) wire n2168_o;
  (* KEEP="TRUE" *) wire n2169_o;
  (* KEEP="TRUE" *) wire n2170_o;
  (* KEEP="TRUE" *) wire n2171_o;
  (* KEEP="TRUE" *) wire n2172_o;
  (* KEEP="TRUE" *) wire n2173_o;
  (* KEEP="TRUE" *) wire n2174_o;
  (* KEEP="TRUE" *) wire n2175_o;
  (* KEEP="TRUE" *) wire n2176_o;
  (* KEEP="TRUE" *) wire n2177_o;
  (* KEEP="TRUE" *) wire n2178_o;
  (* KEEP="TRUE" *) wire n2179_o;
  (* KEEP="TRUE" *) wire n2180_o;
  (* KEEP="TRUE" *) wire n2181_o;
  (* KEEP="TRUE" *) wire n2182_o;
  (* KEEP="TRUE" *) wire n2183_o;
  (* KEEP="TRUE" *) wire n2184_o;
  (* KEEP="TRUE" *) wire n2185_o;
  (* KEEP="TRUE" *) wire n2186_o;
  (* KEEP="TRUE" *) wire n2187_o;
  (* KEEP="TRUE" *) wire n2188_o;
  (* KEEP="TRUE" *) wire n2189_o;
  (* KEEP="TRUE" *) wire n2190_o;
  (* KEEP="TRUE" *) wire n2191_o;
  (* KEEP="TRUE" *) wire n2192_o;
  (* KEEP="TRUE" *) wire n2193_o;
  (* KEEP="TRUE" *) wire n2194_o;
  (* KEEP="TRUE" *) wire n2195_o;
  (* KEEP="TRUE" *) wire n2196_o;
  (* KEEP="TRUE" *) wire n2197_o;
  (* KEEP="TRUE" *) wire n2198_o;
  (* KEEP="TRUE" *) wire n2199_o;
  (* KEEP="TRUE" *) wire n2200_o;
  (* KEEP="TRUE" *) wire n2201_o;
  (* KEEP="TRUE" *) wire n2202_o;
  (* KEEP="TRUE" *) wire n2203_o;
  (* KEEP="TRUE" *) wire n2204_o;
  (* KEEP="TRUE" *) wire n2205_o;
  (* KEEP="TRUE" *) wire n2206_o;
  (* KEEP="TRUE" *) wire n2207_o;
  (* KEEP="TRUE" *) wire n2208_o;
  (* KEEP="TRUE" *) wire n2209_o;
  (* KEEP="TRUE" *) wire n2210_o;
  (* KEEP="TRUE" *) wire n2211_o;
  (* KEEP="TRUE" *) wire n2212_o;
  (* KEEP="TRUE" *) wire n2213_o;
  (* KEEP="TRUE" *) wire n2214_o;
  (* KEEP="TRUE" *) wire n2215_o;
  (* KEEP="TRUE" *) wire n2216_o;
  (* KEEP="TRUE" *) wire n2217_o;
  (* KEEP="TRUE" *) wire n2218_o;
  (* KEEP="TRUE" *) wire n2219_o;
  (* KEEP="TRUE" *) wire n2220_o;
  (* KEEP="TRUE" *) wire n2221_o;
  (* KEEP="TRUE" *) wire n2222_o;
  (* KEEP="TRUE" *) wire n2223_o;
  (* KEEP="TRUE" *) wire n2224_o;
  (* KEEP="TRUE" *) wire n2225_o;
  (* KEEP="TRUE" *) wire n2226_o;
  (* KEEP="TRUE" *) wire n2227_o;
  (* KEEP="TRUE" *) wire n2228_o;
  (* KEEP="TRUE" *) wire n2229_o;
  (* KEEP="TRUE" *) wire n2230_o;
  (* KEEP="TRUE" *) wire n2231_o;
  (* KEEP="TRUE" *) wire n2232_o;
  (* KEEP="TRUE" *) wire n2233_o;
  (* KEEP="TRUE" *) wire n2234_o;
  (* KEEP="TRUE" *) wire n2235_o;
  (* KEEP="TRUE" *) wire n2236_o;
  (* KEEP="TRUE" *) wire n2237_o;
  (* KEEP="TRUE" *) wire n2238_o;
  (* KEEP="TRUE" *) wire n2239_o;
  (* KEEP="TRUE" *) wire n2240_o;
  (* KEEP="TRUE" *) wire n2241_o;
  (* KEEP="TRUE" *) wire n2242_o;
  (* KEEP="TRUE" *) wire n2243_o;
  (* KEEP="TRUE" *) wire n2244_o;
  (* KEEP="TRUE" *) wire n2245_o;
  (* KEEP="TRUE" *) wire n2246_o;
  (* KEEP="TRUE" *) wire n2247_o;
  (* KEEP="TRUE" *) wire n2248_o;
  (* KEEP="TRUE" *) wire n2249_o;
  (* KEEP="TRUE" *) wire n2250_o;
  (* KEEP="TRUE" *) wire n2251_o;
  (* KEEP="TRUE" *) wire n2252_o;
  (* KEEP="TRUE" *) wire n2253_o;
  (* KEEP="TRUE" *) wire n2254_o;
  (* KEEP="TRUE" *) wire n2255_o;
  (* KEEP="TRUE" *) wire n2256_o;
  (* KEEP="TRUE" *) wire n2257_o;
  (* KEEP="TRUE" *) wire n2258_o;
  (* KEEP="TRUE" *) wire n2259_o;
  (* KEEP="TRUE" *) wire n2260_o;
  (* KEEP="TRUE" *) wire n2261_o;
  (* KEEP="TRUE" *) wire n2262_o;
  (* KEEP="TRUE" *) wire n2263_o;
  (* KEEP="TRUE" *) wire n2264_o;
  (* KEEP="TRUE" *) wire n2265_o;
  (* KEEP="TRUE" *) wire n2266_o;
  (* KEEP="TRUE" *) wire n2267_o;
  (* KEEP="TRUE" *) wire n2268_o;
  (* KEEP="TRUE" *) wire n2269_o;
  (* KEEP="TRUE" *) wire n2270_o;
  (* KEEP="TRUE" *) wire n2271_o;
  (* KEEP="TRUE" *) wire n2272_o;
  (* KEEP="TRUE" *) wire n2273_o;
  (* KEEP="TRUE" *) wire n2274_o;
  (* KEEP="TRUE" *) wire n2275_o;
  (* KEEP="TRUE" *) wire n2276_o;
  (* KEEP="TRUE" *) wire n2277_o;
  (* KEEP="TRUE" *) wire n2278_o;
  (* KEEP="TRUE" *) wire n2279_o;
  (* KEEP="TRUE" *) wire n2280_o;
  (* KEEP="TRUE" *) wire n2281_o;
  (* KEEP="TRUE" *) wire n2282_o;
  (* KEEP="TRUE" *) wire n2283_o;
  (* KEEP="TRUE" *) wire n2284_o;
  (* KEEP="TRUE" *) wire n2285_o;
  (* KEEP="TRUE" *) wire n2286_o;
  (* KEEP="TRUE" *) wire n2287_o;
  (* KEEP="TRUE" *) wire n2288_o;
  (* KEEP="TRUE" *) wire n2289_o;
  (* KEEP="TRUE" *) wire n2290_o;
  (* KEEP="TRUE" *) wire n2291_o;
  (* KEEP="TRUE" *) wire n2292_o;
  (* KEEP="TRUE" *) wire n2293_o;
  (* KEEP="TRUE" *) wire n2294_o;
  (* KEEP="TRUE" *) wire n2295_o;
  (* KEEP="TRUE" *) wire n2296_o;
  (* KEEP="TRUE" *) wire n2297_o;
  (* KEEP="TRUE" *) wire n2298_o;
  (* KEEP="TRUE" *) wire n2299_o;
  (* KEEP="TRUE" *) wire n2300_o;
  (* KEEP="TRUE" *) wire n2301_o;
  (* KEEP="TRUE" *) wire n2302_o;
  (* KEEP="TRUE" *) wire n2303_o;
  (* KEEP="TRUE" *) wire n2304_o;
  (* KEEP="TRUE" *) wire n2305_o;
  (* KEEP="TRUE" *) wire n2306_o;
  (* KEEP="TRUE" *) wire n2307_o;
  (* KEEP="TRUE" *) wire n2308_o;
  (* KEEP="TRUE" *) wire n2309_o;
  (* KEEP="TRUE" *) wire n2310_o;
  (* KEEP="TRUE" *) wire n2311_o;
  (* KEEP="TRUE" *) wire n2312_o;
  (* KEEP="TRUE" *) wire n2313_o;
  (* KEEP="TRUE" *) wire n2314_o;
  (* KEEP="TRUE" *) wire n2315_o;
  (* KEEP="TRUE" *) wire n2316_o;
  (* KEEP="TRUE" *) wire n2317_o;
  (* KEEP="TRUE" *) wire n2318_o;
  (* KEEP="TRUE" *) wire n2319_o;
  (* KEEP="TRUE" *) wire n2320_o;
  (* KEEP="TRUE" *) wire n2321_o;
  (* KEEP="TRUE" *) wire n2322_o;
  (* KEEP="TRUE" *) wire n2323_o;
  (* KEEP="TRUE" *) wire n2324_o;
  (* KEEP="TRUE" *) wire n2325_o;
  (* KEEP="TRUE" *) wire n2326_o;
  (* KEEP="TRUE" *) wire n2327_o;
  (* KEEP="TRUE" *) wire n2328_o;
  (* KEEP="TRUE" *) wire n2329_o;
  (* KEEP="TRUE" *) wire n2330_o;
  (* KEEP="TRUE" *) wire n2331_o;
  (* KEEP="TRUE" *) wire n2332_o;
  (* KEEP="TRUE" *) wire n2333_o;
  (* KEEP="TRUE" *) wire n2334_o;
  (* KEEP="TRUE" *) wire n2335_o;
  (* KEEP="TRUE" *) wire n2336_o;
  (* KEEP="TRUE" *) wire n2337_o;
  (* KEEP="TRUE" *) wire n2338_o;
  (* KEEP="TRUE" *) wire n2339_o;
  (* KEEP="TRUE" *) wire n2340_o;
  (* KEEP="TRUE" *) wire n2341_o;
  (* KEEP="TRUE" *) wire n2342_o;
  (* KEEP="TRUE" *) wire n2343_o;
  (* KEEP="TRUE" *) wire n2344_o;
  (* KEEP="TRUE" *) wire n2345_o;
  (* KEEP="TRUE" *) wire n2346_o;
  (* KEEP="TRUE" *) wire n2347_o;
  (* KEEP="TRUE" *) wire n2348_o;
  (* KEEP="TRUE" *) wire n2349_o;
  (* KEEP="TRUE" *) wire n2350_o;
  (* KEEP="TRUE" *) wire n2351_o;
  (* KEEP="TRUE" *) wire n2352_o;
  (* KEEP="TRUE" *) wire n2353_o;
  (* KEEP="TRUE" *) wire n2354_o;
  (* KEEP="TRUE" *) wire n2355_o;
  (* KEEP="TRUE" *) wire n2356_o;
  (* KEEP="TRUE" *) wire n2357_o;
  (* KEEP="TRUE" *) wire n2358_o;
  (* KEEP="TRUE" *) wire n2359_o;
  (* KEEP="TRUE" *) wire n2360_o;
  (* KEEP="TRUE" *) wire n2361_o;
  (* KEEP="TRUE" *) wire n2362_o;
  (* KEEP="TRUE" *) wire n2363_o;
  (* KEEP="TRUE" *) wire n2364_o;
  (* KEEP="TRUE" *) wire n2365_o;
  (* KEEP="TRUE" *) wire n2366_o;
  (* KEEP="TRUE" *) wire n2367_o;
  (* KEEP="TRUE" *) wire n2368_o;
  (* KEEP="TRUE" *) wire n2369_o;
  (* KEEP="TRUE" *) wire n2370_o;
  (* KEEP="TRUE" *) wire n2371_o;
  (* KEEP="TRUE" *) wire n2372_o;
  (* KEEP="TRUE" *) wire n2373_o;
  (* KEEP="TRUE" *) wire n2374_o;
  (* KEEP="TRUE" *) wire n2375_o;
  (* KEEP="TRUE" *) wire n2376_o;
  (* KEEP="TRUE" *) wire n2377_o;
  (* KEEP="TRUE" *) wire n2378_o;
  (* KEEP="TRUE" *) wire n2379_o;
  (* KEEP="TRUE" *) wire n2380_o;
  (* KEEP="TRUE" *) wire n2381_o;
  (* KEEP="TRUE" *) wire n2382_o;
  (* KEEP="TRUE" *) wire n2383_o;
  (* KEEP="TRUE" *) wire n2384_o;
  (* KEEP="TRUE" *) wire n2385_o;
  (* KEEP="TRUE" *) wire n2386_o;
  (* KEEP="TRUE" *) wire n2387_o;
  (* KEEP="TRUE" *) wire n2388_o;
  (* KEEP="TRUE" *) wire n2389_o;
  (* KEEP="TRUE" *) wire n2390_o;
  (* KEEP="TRUE" *) wire n2391_o;
  (* KEEP="TRUE" *) wire n2392_o;
  (* KEEP="TRUE" *) wire n2393_o;
  (* KEEP="TRUE" *) wire n2394_o;
  (* KEEP="TRUE" *) wire n2395_o;
  (* KEEP="TRUE" *) wire n2396_o;
  (* KEEP="TRUE" *) wire n2397_o;
  (* KEEP="TRUE" *) wire n2398_o;
  (* KEEP="TRUE" *) wire n2399_o;
  (* KEEP="TRUE" *) wire n2400_o;
  (* KEEP="TRUE" *) wire n2401_o;
  (* KEEP="TRUE" *) wire n2402_o;
  (* KEEP="TRUE" *) wire n2403_o;
  (* KEEP="TRUE" *) wire n2404_o;
  (* KEEP="TRUE" *) wire n2405_o;
  (* KEEP="TRUE" *) wire n2406_o;
  (* KEEP="TRUE" *) wire n2407_o;
  (* KEEP="TRUE" *) wire n2408_o;
  (* KEEP="TRUE" *) wire n2409_o;
  (* KEEP="TRUE" *) wire n2410_o;
  (* KEEP="TRUE" *) wire n2411_o;
  (* KEEP="TRUE" *) wire n2412_o;
  (* KEEP="TRUE" *) wire n2413_o;
  (* KEEP="TRUE" *) wire n2414_o;
  (* KEEP="TRUE" *) wire n2415_o;
  (* KEEP="TRUE" *) wire n2416_o;
  (* KEEP="TRUE" *) wire n2417_o;
  (* KEEP="TRUE" *) wire n2418_o;
  (* KEEP="TRUE" *) wire n2419_o;
  (* KEEP="TRUE" *) wire n2420_o;
  (* KEEP="TRUE" *) wire n2421_o;
  (* KEEP="TRUE" *) wire n2422_o;
  (* KEEP="TRUE" *) wire n2423_o;
  (* KEEP="TRUE" *) wire n2424_o;
  (* KEEP="TRUE" *) wire n2425_o;
  (* KEEP="TRUE" *) wire n2426_o;
  (* KEEP="TRUE" *) wire n2427_o;
  (* KEEP="TRUE" *) wire n2428_o;
  (* KEEP="TRUE" *) wire n2429_o;
  (* KEEP="TRUE" *) wire n2430_o;
  (* KEEP="TRUE" *) wire n2431_o;
  (* KEEP="TRUE" *) wire n2432_o;
  (* KEEP="TRUE" *) wire n2433_o;
  (* KEEP="TRUE" *) wire n2434_o;
  (* KEEP="TRUE" *) wire n2435_o;
  (* KEEP="TRUE" *) wire n2436_o;
  (* KEEP="TRUE" *) wire n2437_o;
  (* KEEP="TRUE" *) wire n2438_o;
  (* KEEP="TRUE" *) wire n2439_o;
  (* KEEP="TRUE" *) wire n2440_o;
  (* KEEP="TRUE" *) wire n2441_o;
  (* KEEP="TRUE" *) wire n2442_o;
  (* KEEP="TRUE" *) wire n2443_o;
  (* KEEP="TRUE" *) wire n2444_o;
  (* KEEP="TRUE" *) wire n2445_o;
  (* KEEP="TRUE" *) wire n2446_o;
  (* KEEP="TRUE" *) wire n2447_o;
  (* KEEP="TRUE" *) wire n2448_o;
  (* KEEP="TRUE" *) wire n2449_o;
  (* KEEP="TRUE" *) wire n2450_o;
  (* KEEP="TRUE" *) wire n2451_o;
  (* KEEP="TRUE" *) wire n2452_o;
  (* KEEP="TRUE" *) wire n2453_o;
  (* KEEP="TRUE" *) wire n2454_o;
  (* KEEP="TRUE" *) wire n2455_o;
  (* KEEP="TRUE" *) wire n2456_o;
  (* KEEP="TRUE" *) wire n2457_o;
  (* KEEP="TRUE" *) wire n2458_o;
  (* KEEP="TRUE" *) wire n2459_o;
  (* KEEP="TRUE" *) wire n2460_o;
  (* KEEP="TRUE" *) wire n2461_o;
  (* KEEP="TRUE" *) wire n2462_o;
  (* KEEP="TRUE" *) wire n2463_o;
  (* KEEP="TRUE" *) wire n2464_o;
  (* KEEP="TRUE" *) wire n2465_o;
  (* KEEP="TRUE" *) wire n2466_o;
  (* KEEP="TRUE" *) wire n2467_o;
  (* KEEP="TRUE" *) wire n2468_o;
  (* KEEP="TRUE" *) wire n2469_o;
  (* KEEP="TRUE" *) wire n2470_o;
  (* KEEP="TRUE" *) wire n2471_o;
  (* KEEP="TRUE" *) wire n2472_o;
  (* KEEP="TRUE" *) wire n2473_o;
  (* KEEP="TRUE" *) wire n2474_o;
  (* KEEP="TRUE" *) wire n2475_o;
  (* KEEP="TRUE" *) wire n2476_o;
  (* KEEP="TRUE" *) wire n2477_o;
  (* KEEP="TRUE" *) wire n2478_o;
  (* KEEP="TRUE" *) wire n2479_o;
  (* KEEP="TRUE" *) wire n2480_o;
  (* KEEP="TRUE" *) wire n2481_o;
  (* KEEP="TRUE" *) wire n2482_o;
  (* KEEP="TRUE" *) wire n2483_o;
  (* KEEP="TRUE" *) wire n2484_o;
  (* KEEP="TRUE" *) wire n2485_o;
  (* KEEP="TRUE" *) wire n2486_o;
  (* KEEP="TRUE" *) wire n2487_o;
  (* KEEP="TRUE" *) wire n2488_o;
  (* KEEP="TRUE" *) wire n2489_o;
  (* KEEP="TRUE" *) wire n2490_o;
  (* KEEP="TRUE" *) wire n2491_o;
  (* KEEP="TRUE" *) wire n2492_o;
  (* KEEP="TRUE" *) wire n2493_o;
  (* KEEP="TRUE" *) wire n2494_o;
  (* KEEP="TRUE" *) wire n2495_o;
  (* KEEP="TRUE" *) wire n2496_o;
  (* KEEP="TRUE" *) wire n2497_o;
  (* KEEP="TRUE" *) wire n2498_o;
  (* KEEP="TRUE" *) wire n2499_o;
  (* KEEP="TRUE" *) wire n2500_o;
  (* KEEP="TRUE" *) wire n2501_o;
  (* KEEP="TRUE" *) wire n2502_o;
  (* KEEP="TRUE" *) wire n2503_o;
  (* KEEP="TRUE" *) wire n2504_o;
  (* KEEP="TRUE" *) wire n2505_o;
  (* KEEP="TRUE" *) wire n2506_o;
  (* KEEP="TRUE" *) wire n2507_o;
  (* KEEP="TRUE" *) wire n2508_o;
  (* KEEP="TRUE" *) wire n2509_o;
  (* KEEP="TRUE" *) wire n2510_o;
  (* KEEP="TRUE" *) wire n2511_o;
  (* KEEP="TRUE" *) wire n2512_o;
  (* KEEP="TRUE" *) wire n2513_o;
  (* KEEP="TRUE" *) wire n2514_o;
  (* KEEP="TRUE" *) wire n2515_o;
  (* KEEP="TRUE" *) wire n2516_o;
  (* KEEP="TRUE" *) wire n2517_o;
  (* KEEP="TRUE" *) wire n2518_o;
  (* KEEP="TRUE" *) wire n2519_o;
  (* KEEP="TRUE" *) wire n2520_o;
  (* KEEP="TRUE" *) wire n2521_o;
  (* KEEP="TRUE" *) wire n2522_o;
  (* KEEP="TRUE" *) wire n2523_o;
  (* KEEP="TRUE" *) wire n2524_o;
  (* KEEP="TRUE" *) wire n2525_o;
  (* KEEP="TRUE" *) wire n2526_o;
  (* KEEP="TRUE" *) wire n2527_o;
  (* KEEP="TRUE" *) wire n2528_o;
  (* KEEP="TRUE" *) wire n2529_o;
  (* KEEP="TRUE" *) wire n2530_o;
  (* KEEP="TRUE" *) wire n2531_o;
  (* KEEP="TRUE" *) wire n2532_o;
  (* KEEP="TRUE" *) wire n2533_o;
  (* KEEP="TRUE" *) wire n2534_o;
  (* KEEP="TRUE" *) wire n2535_o;
  (* KEEP="TRUE" *) wire n2536_o;
  (* KEEP="TRUE" *) wire n2537_o;
  (* KEEP="TRUE" *) wire n2538_o;
  (* KEEP="TRUE" *) wire n2539_o;
  (* KEEP="TRUE" *) wire n2540_o;
  (* KEEP="TRUE" *) wire n2541_o;
  (* KEEP="TRUE" *) wire n2542_o;
  (* KEEP="TRUE" *) wire n2543_o;
  (* KEEP="TRUE" *) wire n2544_o;
  (* KEEP="TRUE" *) wire n2545_o;
  (* KEEP="TRUE" *) wire n2546_o;
  (* KEEP="TRUE" *) wire n2547_o;
  (* KEEP="TRUE" *) wire n2548_o;
  (* KEEP="TRUE" *) wire n2549_o;
  (* KEEP="TRUE" *) wire n2550_o;
  (* KEEP="TRUE" *) wire n2551_o;
  (* KEEP="TRUE" *) wire n2552_o;
  (* KEEP="TRUE" *) wire n2553_o;
  (* KEEP="TRUE" *) wire n2554_o;
  (* KEEP="TRUE" *) wire n2555_o;
  (* KEEP="TRUE" *) wire n2556_o;
  (* KEEP="TRUE" *) wire n2557_o;
  (* KEEP="TRUE" *) wire n2558_o;
  (* KEEP="TRUE" *) wire n2559_o;
  (* KEEP="TRUE" *) wire n2560_o;
  (* KEEP="TRUE" *) wire n2561_o;
  (* KEEP="TRUE" *) wire n2562_o;
  (* KEEP="TRUE" *) wire n2563_o;
  (* KEEP="TRUE" *) wire n2564_o;
  (* KEEP="TRUE" *) wire n2565_o;
  (* KEEP="TRUE" *) wire n2566_o;
  (* KEEP="TRUE" *) wire n2567_o;
  (* KEEP="TRUE" *) wire n2568_o;
  (* KEEP="TRUE" *) wire n2569_o;
  (* KEEP="TRUE" *) wire [255:0] n2570_o;
  (* KEEP="TRUE" *) wire n2571_o;
  (* KEEP="TRUE" *) wire n2572_o;
  (* KEEP="TRUE" *) wire n2573_o;
  (* KEEP="TRUE" *) wire n2574_o;
  (* KEEP="TRUE" *) wire n2575_o;
  (* KEEP="TRUE" *) wire n2576_o;
  (* KEEP="TRUE" *) wire n2577_o;
  (* KEEP="TRUE" *) wire n2578_o;
  (* KEEP="TRUE" *) wire n2579_o;
  (* KEEP="TRUE" *) wire n2580_o;
  (* KEEP="TRUE" *) wire n2581_o;
  (* KEEP="TRUE" *) wire n2582_o;
  (* KEEP="TRUE" *) wire n2583_o;
  (* KEEP="TRUE" *) wire n2584_o;
  (* KEEP="TRUE" *) wire n2585_o;
  (* KEEP="TRUE" *) wire n2586_o;
  (* KEEP="TRUE" *) wire n2587_o;
  (* KEEP="TRUE" *) wire n2588_o;
  (* KEEP="TRUE" *) wire n2589_o;
  (* KEEP="TRUE" *) wire n2590_o;
  (* KEEP="TRUE" *) wire n2591_o;
  (* KEEP="TRUE" *) wire n2592_o;
  (* KEEP="TRUE" *) wire n2593_o;
  (* KEEP="TRUE" *) wire n2594_o;
  (* KEEP="TRUE" *) wire n2595_o;
  (* KEEP="TRUE" *) wire n2596_o;
  (* KEEP="TRUE" *) wire n2597_o;
  (* KEEP="TRUE" *) wire n2598_o;
  (* KEEP="TRUE" *) wire n2599_o;
  (* KEEP="TRUE" *) wire n2600_o;
  (* KEEP="TRUE" *) wire n2601_o;
  (* KEEP="TRUE" *) wire n2602_o;
  (* KEEP="TRUE" *) wire n2603_o;
  (* KEEP="TRUE" *) wire n2604_o;
  (* KEEP="TRUE" *) wire n2605_o;
  (* KEEP="TRUE" *) wire n2606_o;
  (* KEEP="TRUE" *) wire n2607_o;
  (* KEEP="TRUE" *) wire n2608_o;
  (* KEEP="TRUE" *) wire n2609_o;
  (* KEEP="TRUE" *) wire n2610_o;
  (* KEEP="TRUE" *) wire n2611_o;
  (* KEEP="TRUE" *) wire n2612_o;
  (* KEEP="TRUE" *) wire n2613_o;
  (* KEEP="TRUE" *) wire n2614_o;
  (* KEEP="TRUE" *) wire n2615_o;
  (* KEEP="TRUE" *) wire n2616_o;
  (* KEEP="TRUE" *) wire n2617_o;
  (* KEEP="TRUE" *) wire n2618_o;
  (* KEEP="TRUE" *) wire n2619_o;
  (* KEEP="TRUE" *) wire n2620_o;
  (* KEEP="TRUE" *) wire n2621_o;
  (* KEEP="TRUE" *) wire n2622_o;
  (* KEEP="TRUE" *) wire n2623_o;
  (* KEEP="TRUE" *) wire n2624_o;
  (* KEEP="TRUE" *) wire n2625_o;
  (* KEEP="TRUE" *) wire n2626_o;
  (* KEEP="TRUE" *) wire n2627_o;
  (* KEEP="TRUE" *) wire n2628_o;
  (* KEEP="TRUE" *) wire n2629_o;
  (* KEEP="TRUE" *) wire n2630_o;
  (* KEEP="TRUE" *) wire n2631_o;
  (* KEEP="TRUE" *) wire n2632_o;
  (* KEEP="TRUE" *) wire n2633_o;
  (* KEEP="TRUE" *) wire n2634_o;
  (* KEEP="TRUE" *) wire n2635_o;
  (* KEEP="TRUE" *) wire n2636_o;
  (* KEEP="TRUE" *) wire n2637_o;
  (* KEEP="TRUE" *) wire n2638_o;
  (* KEEP="TRUE" *) wire n2639_o;
  (* KEEP="TRUE" *) wire n2640_o;
  (* KEEP="TRUE" *) wire n2641_o;
  (* KEEP="TRUE" *) wire n2642_o;
  (* KEEP="TRUE" *) wire n2643_o;
  (* KEEP="TRUE" *) wire n2644_o;
  (* KEEP="TRUE" *) wire n2645_o;
  (* KEEP="TRUE" *) wire n2646_o;
  (* KEEP="TRUE" *) wire n2647_o;
  (* KEEP="TRUE" *) wire n2648_o;
  (* KEEP="TRUE" *) wire n2649_o;
  (* KEEP="TRUE" *) wire n2650_o;
  (* KEEP="TRUE" *) wire n2651_o;
  (* KEEP="TRUE" *) wire n2652_o;
  (* KEEP="TRUE" *) wire n2653_o;
  (* KEEP="TRUE" *) wire n2654_o;
  (* KEEP="TRUE" *) wire n2655_o;
  (* KEEP="TRUE" *) wire n2656_o;
  (* KEEP="TRUE" *) wire n2657_o;
  (* KEEP="TRUE" *) wire n2658_o;
  (* KEEP="TRUE" *) wire n2659_o;
  (* KEEP="TRUE" *) wire n2660_o;
  (* KEEP="TRUE" *) wire n2661_o;
  (* KEEP="TRUE" *) wire n2662_o;
  (* KEEP="TRUE" *) wire n2663_o;
  (* KEEP="TRUE" *) wire n2664_o;
  (* KEEP="TRUE" *) wire n2665_o;
  (* KEEP="TRUE" *) wire n2666_o;
  (* KEEP="TRUE" *) wire n2667_o;
  (* KEEP="TRUE" *) wire n2668_o;
  (* KEEP="TRUE" *) wire n2669_o;
  (* KEEP="TRUE" *) wire n2670_o;
  (* KEEP="TRUE" *) wire n2671_o;
  (* KEEP="TRUE" *) wire n2672_o;
  (* KEEP="TRUE" *) wire n2673_o;
  (* KEEP="TRUE" *) wire n2674_o;
  (* KEEP="TRUE" *) wire n2675_o;
  (* KEEP="TRUE" *) wire n2676_o;
  (* KEEP="TRUE" *) wire n2677_o;
  (* KEEP="TRUE" *) wire n2678_o;
  (* KEEP="TRUE" *) wire n2679_o;
  (* KEEP="TRUE" *) wire n2680_o;
  (* KEEP="TRUE" *) wire n2681_o;
  (* KEEP="TRUE" *) wire n2682_o;
  (* KEEP="TRUE" *) wire n2683_o;
  (* KEEP="TRUE" *) wire n2684_o;
  (* KEEP="TRUE" *) wire n2685_o;
  (* KEEP="TRUE" *) wire n2686_o;
  (* KEEP="TRUE" *) wire n2687_o;
  (* KEEP="TRUE" *) wire n2688_o;
  (* KEEP="TRUE" *) wire n2689_o;
  (* KEEP="TRUE" *) wire n2690_o;
  (* KEEP="TRUE" *) wire n2691_o;
  (* KEEP="TRUE" *) wire n2692_o;
  (* KEEP="TRUE" *) wire n2693_o;
  (* KEEP="TRUE" *) wire n2694_o;
  (* KEEP="TRUE" *) wire n2695_o;
  (* KEEP="TRUE" *) wire n2696_o;
  (* KEEP="TRUE" *) wire n2697_o;
  (* KEEP="TRUE" *) wire n2698_o;
  (* KEEP="TRUE" *) wire n2699_o;
  (* KEEP="TRUE" *) wire n2700_o;
  (* KEEP="TRUE" *) wire n2701_o;
  (* KEEP="TRUE" *) wire n2702_o;
  (* KEEP="TRUE" *) wire n2703_o;
  (* KEEP="TRUE" *) wire n2704_o;
  (* KEEP="TRUE" *) wire n2705_o;
  (* KEEP="TRUE" *) wire n2706_o;
  (* KEEP="TRUE" *) wire n2707_o;
  (* KEEP="TRUE" *) wire n2708_o;
  (* KEEP="TRUE" *) wire n2709_o;
  (* KEEP="TRUE" *) wire n2710_o;
  (* KEEP="TRUE" *) wire n2711_o;
  (* KEEP="TRUE" *) wire n2712_o;
  (* KEEP="TRUE" *) wire n2713_o;
  (* KEEP="TRUE" *) wire n2714_o;
  (* KEEP="TRUE" *) wire n2715_o;
  (* KEEP="TRUE" *) wire n2716_o;
  (* KEEP="TRUE" *) wire n2717_o;
  (* KEEP="TRUE" *) wire n2718_o;
  (* KEEP="TRUE" *) wire n2719_o;
  (* KEEP="TRUE" *) wire n2720_o;
  (* KEEP="TRUE" *) wire n2721_o;
  (* KEEP="TRUE" *) wire n2722_o;
  (* KEEP="TRUE" *) wire n2723_o;
  (* KEEP="TRUE" *) wire n2724_o;
  (* KEEP="TRUE" *) wire n2725_o;
  (* KEEP="TRUE" *) wire n2726_o;
  (* KEEP="TRUE" *) wire n2727_o;
  (* KEEP="TRUE" *) wire n2728_o;
  (* KEEP="TRUE" *) wire n2729_o;
  (* KEEP="TRUE" *) wire n2730_o;
  (* KEEP="TRUE" *) wire n2731_o;
  (* KEEP="TRUE" *) wire n2732_o;
  (* KEEP="TRUE" *) wire n2733_o;
  (* KEEP="TRUE" *) wire n2734_o;
  (* KEEP="TRUE" *) wire n2735_o;
  (* KEEP="TRUE" *) wire n2736_o;
  (* KEEP="TRUE" *) wire n2737_o;
  (* KEEP="TRUE" *) wire n2738_o;
  (* KEEP="TRUE" *) wire n2739_o;
  (* KEEP="TRUE" *) wire n2740_o;
  (* KEEP="TRUE" *) wire n2741_o;
  (* KEEP="TRUE" *) wire n2742_o;
  (* KEEP="TRUE" *) wire n2743_o;
  (* KEEP="TRUE" *) wire n2744_o;
  (* KEEP="TRUE" *) wire n2745_o;
  (* KEEP="TRUE" *) wire n2746_o;
  (* KEEP="TRUE" *) wire n2747_o;
  (* KEEP="TRUE" *) wire n2748_o;
  (* KEEP="TRUE" *) wire n2749_o;
  (* KEEP="TRUE" *) wire n2750_o;
  (* KEEP="TRUE" *) wire n2751_o;
  (* KEEP="TRUE" *) wire n2752_o;
  (* KEEP="TRUE" *) wire n2753_o;
  (* KEEP="TRUE" *) wire n2754_o;
  (* KEEP="TRUE" *) wire n2755_o;
  (* KEEP="TRUE" *) wire n2756_o;
  (* KEEP="TRUE" *) wire n2757_o;
  (* KEEP="TRUE" *) wire n2758_o;
  (* KEEP="TRUE" *) wire n2759_o;
  (* KEEP="TRUE" *) wire n2760_o;
  (* KEEP="TRUE" *) wire n2761_o;
  (* KEEP="TRUE" *) wire n2762_o;
  (* KEEP="TRUE" *) wire n2763_o;
  (* KEEP="TRUE" *) wire n2764_o;
  (* KEEP="TRUE" *) wire n2765_o;
  (* KEEP="TRUE" *) wire n2766_o;
  (* KEEP="TRUE" *) wire n2767_o;
  (* KEEP="TRUE" *) wire n2768_o;
  (* KEEP="TRUE" *) wire n2769_o;
  (* KEEP="TRUE" *) wire n2770_o;
  (* KEEP="TRUE" *) wire n2771_o;
  (* KEEP="TRUE" *) wire n2772_o;
  (* KEEP="TRUE" *) wire n2773_o;
  (* KEEP="TRUE" *) wire n2774_o;
  (* KEEP="TRUE" *) wire n2775_o;
  (* KEEP="TRUE" *) wire n2776_o;
  (* KEEP="TRUE" *) wire n2777_o;
  (* KEEP="TRUE" *) wire n2778_o;
  (* KEEP="TRUE" *) wire n2779_o;
  (* KEEP="TRUE" *) wire n2780_o;
  (* KEEP="TRUE" *) wire n2781_o;
  (* KEEP="TRUE" *) wire n2782_o;
  (* KEEP="TRUE" *) wire n2783_o;
  (* KEEP="TRUE" *) wire n2784_o;
  (* KEEP="TRUE" *) wire n2785_o;
  (* KEEP="TRUE" *) wire n2786_o;
  (* KEEP="TRUE" *) wire n2787_o;
  (* KEEP="TRUE" *) wire n2788_o;
  (* KEEP="TRUE" *) wire n2789_o;
  (* KEEP="TRUE" *) wire n2790_o;
  (* KEEP="TRUE" *) wire n2791_o;
  (* KEEP="TRUE" *) wire n2792_o;
  (* KEEP="TRUE" *) wire n2793_o;
  (* KEEP="TRUE" *) wire n2794_o;
  (* KEEP="TRUE" *) wire n2795_o;
  (* KEEP="TRUE" *) wire n2796_o;
  (* KEEP="TRUE" *) wire n2797_o;
  (* KEEP="TRUE" *) wire n2798_o;
  (* KEEP="TRUE" *) wire n2799_o;
  (* KEEP="TRUE" *) wire n2800_o;
  (* KEEP="TRUE" *) wire n2801_o;
  (* KEEP="TRUE" *) wire n2802_o;
  (* KEEP="TRUE" *) wire n2803_o;
  (* KEEP="TRUE" *) wire n2804_o;
  (* KEEP="TRUE" *) wire n2805_o;
  (* KEEP="TRUE" *) wire n2806_o;
  (* KEEP="TRUE" *) wire n2807_o;
  (* KEEP="TRUE" *) wire n2808_o;
  (* KEEP="TRUE" *) wire n2809_o;
  (* KEEP="TRUE" *) wire n2810_o;
  (* KEEP="TRUE" *) wire n2811_o;
  (* KEEP="TRUE" *) wire n2812_o;
  (* KEEP="TRUE" *) wire n2813_o;
  (* KEEP="TRUE" *) wire n2814_o;
  (* KEEP="TRUE" *) wire n2815_o;
  (* KEEP="TRUE" *) wire n2816_o;
  (* KEEP="TRUE" *) wire n2817_o;
  (* KEEP="TRUE" *) wire n2818_o;
  (* KEEP="TRUE" *) wire n2819_o;
  (* KEEP="TRUE" *) wire n2820_o;
  (* KEEP="TRUE" *) wire n2821_o;
  (* KEEP="TRUE" *) wire n2822_o;
  (* KEEP="TRUE" *) wire n2823_o;
  (* KEEP="TRUE" *) wire n2824_o;
  (* KEEP="TRUE" *) wire n2825_o;
  (* KEEP="TRUE" *) wire n2826_o;
  (* KEEP="TRUE" *) wire n2827_o;
  (* KEEP="TRUE" *) wire n2828_o;
  (* KEEP="TRUE" *) wire n2829_o;
  (* KEEP="TRUE" *) wire n2830_o;
  (* KEEP="TRUE" *) wire n2831_o;
  (* KEEP="TRUE" *) wire n2832_o;
  (* KEEP="TRUE" *) wire n2833_o;
  (* KEEP="TRUE" *) wire n2834_o;
  (* KEEP="TRUE" *) wire n2835_o;
  (* KEEP="TRUE" *) wire n2836_o;
  (* KEEP="TRUE" *) wire n2837_o;
  (* KEEP="TRUE" *) wire n2838_o;
  (* KEEP="TRUE" *) wire n2839_o;
  (* KEEP="TRUE" *) wire n2840_o;
  (* KEEP="TRUE" *) wire n2841_o;
  (* KEEP="TRUE" *) wire n2842_o;
  (* KEEP="TRUE" *) wire n2843_o;
  (* KEEP="TRUE" *) wire n2844_o;
  (* KEEP="TRUE" *) wire n2845_o;
  (* KEEP="TRUE" *) wire n2846_o;
  (* KEEP="TRUE" *) wire n2847_o;
  (* KEEP="TRUE" *) wire n2848_o;
  (* KEEP="TRUE" *) wire n2849_o;
  (* KEEP="TRUE" *) wire n2850_o;
  (* KEEP="TRUE" *) wire n2851_o;
  (* KEEP="TRUE" *) wire n2852_o;
  (* KEEP="TRUE" *) wire n2853_o;
  (* KEEP="TRUE" *) wire n2854_o;
  (* KEEP="TRUE" *) wire n2855_o;
  (* KEEP="TRUE" *) wire n2856_o;
  (* KEEP="TRUE" *) wire n2857_o;
  (* KEEP="TRUE" *) wire n2858_o;
  (* KEEP="TRUE" *) wire n2859_o;
  (* KEEP="TRUE" *) wire n2860_o;
  (* KEEP="TRUE" *) wire n2861_o;
  (* KEEP="TRUE" *) wire n2862_o;
  (* KEEP="TRUE" *) wire n2863_o;
  (* KEEP="TRUE" *) wire n2864_o;
  (* KEEP="TRUE" *) wire n2865_o;
  (* KEEP="TRUE" *) wire n2866_o;
  (* KEEP="TRUE" *) wire n2867_o;
  (* KEEP="TRUE" *) wire n2868_o;
  (* KEEP="TRUE" *) wire n2869_o;
  (* KEEP="TRUE" *) wire n2870_o;
  (* KEEP="TRUE" *) wire n2871_o;
  (* KEEP="TRUE" *) wire n2872_o;
  (* KEEP="TRUE" *) wire n2873_o;
  (* KEEP="TRUE" *) wire n2874_o;
  (* KEEP="TRUE" *) wire n2875_o;
  (* KEEP="TRUE" *) wire n2876_o;
  (* KEEP="TRUE" *) wire n2877_o;
  (* KEEP="TRUE" *) wire n2878_o;
  (* KEEP="TRUE" *) wire n2879_o;
  (* KEEP="TRUE" *) wire n2880_o;
  (* KEEP="TRUE" *) wire n2881_o;
  (* KEEP="TRUE" *) wire n2882_o;
  (* KEEP="TRUE" *) wire n2883_o;
  (* KEEP="TRUE" *) wire n2884_o;
  (* KEEP="TRUE" *) wire n2885_o;
  (* KEEP="TRUE" *) wire n2886_o;
  (* KEEP="TRUE" *) wire n2887_o;
  (* KEEP="TRUE" *) wire n2888_o;
  (* KEEP="TRUE" *) wire n2889_o;
  (* KEEP="TRUE" *) wire n2890_o;
  (* KEEP="TRUE" *) wire n2891_o;
  (* KEEP="TRUE" *) wire n2892_o;
  (* KEEP="TRUE" *) wire n2893_o;
  (* KEEP="TRUE" *) wire n2894_o;
  (* KEEP="TRUE" *) wire n2895_o;
  (* KEEP="TRUE" *) wire n2896_o;
  (* KEEP="TRUE" *) wire n2897_o;
  (* KEEP="TRUE" *) wire n2898_o;
  (* KEEP="TRUE" *) wire n2899_o;
  (* KEEP="TRUE" *) wire n2900_o;
  (* KEEP="TRUE" *) wire n2901_o;
  (* KEEP="TRUE" *) wire n2902_o;
  (* KEEP="TRUE" *) wire n2903_o;
  (* KEEP="TRUE" *) wire n2904_o;
  (* KEEP="TRUE" *) wire n2905_o;
  (* KEEP="TRUE" *) wire n2906_o;
  (* KEEP="TRUE" *) wire n2907_o;
  (* KEEP="TRUE" *) wire n2908_o;
  (* KEEP="TRUE" *) wire n2909_o;
  (* KEEP="TRUE" *) wire n2910_o;
  (* KEEP="TRUE" *) wire n2911_o;
  (* KEEP="TRUE" *) wire n2912_o;
  (* KEEP="TRUE" *) wire n2913_o;
  (* KEEP="TRUE" *) wire n2914_o;
  (* KEEP="TRUE" *) wire n2915_o;
  (* KEEP="TRUE" *) wire n2916_o;
  (* KEEP="TRUE" *) wire n2917_o;
  (* KEEP="TRUE" *) wire n2918_o;
  (* KEEP="TRUE" *) wire n2919_o;
  (* KEEP="TRUE" *) wire n2920_o;
  (* KEEP="TRUE" *) wire n2921_o;
  (* KEEP="TRUE" *) wire n2922_o;
  (* KEEP="TRUE" *) wire n2923_o;
  (* KEEP="TRUE" *) wire n2924_o;
  (* KEEP="TRUE" *) wire n2925_o;
  (* KEEP="TRUE" *) wire n2926_o;
  (* KEEP="TRUE" *) wire n2927_o;
  (* KEEP="TRUE" *) wire n2928_o;
  (* KEEP="TRUE" *) wire n2929_o;
  (* KEEP="TRUE" *) wire n2930_o;
  (* KEEP="TRUE" *) wire n2931_o;
  (* KEEP="TRUE" *) wire n2932_o;
  (* KEEP="TRUE" *) wire n2933_o;
  (* KEEP="TRUE" *) wire n2934_o;
  (* KEEP="TRUE" *) wire n2935_o;
  (* KEEP="TRUE" *) wire n2936_o;
  (* KEEP="TRUE" *) wire n2937_o;
  (* KEEP="TRUE" *) wire n2938_o;
  (* KEEP="TRUE" *) wire n2939_o;
  (* KEEP="TRUE" *) wire n2940_o;
  (* KEEP="TRUE" *) wire n2941_o;
  (* KEEP="TRUE" *) wire n2942_o;
  (* KEEP="TRUE" *) wire n2943_o;
  (* KEEP="TRUE" *) wire n2944_o;
  (* KEEP="TRUE" *) wire n2945_o;
  (* KEEP="TRUE" *) wire n2946_o;
  (* KEEP="TRUE" *) wire n2947_o;
  (* KEEP="TRUE" *) wire n2948_o;
  (* KEEP="TRUE" *) wire n2949_o;
  (* KEEP="TRUE" *) wire n2950_o;
  (* KEEP="TRUE" *) wire n2951_o;
  (* KEEP="TRUE" *) wire n2952_o;
  (* KEEP="TRUE" *) wire n2953_o;
  (* KEEP="TRUE" *) wire n2954_o;
  (* KEEP="TRUE" *) wire n2955_o;
  (* KEEP="TRUE" *) wire n2956_o;
  (* KEEP="TRUE" *) wire n2957_o;
  (* KEEP="TRUE" *) wire n2958_o;
  (* KEEP="TRUE" *) wire n2959_o;
  (* KEEP="TRUE" *) wire n2960_o;
  (* KEEP="TRUE" *) wire n2961_o;
  (* KEEP="TRUE" *) wire n2962_o;
  (* KEEP="TRUE" *) wire n2963_o;
  (* KEEP="TRUE" *) wire n2964_o;
  (* KEEP="TRUE" *) wire n2965_o;
  (* KEEP="TRUE" *) wire n2966_o;
  (* KEEP="TRUE" *) wire n2967_o;
  (* KEEP="TRUE" *) wire n2968_o;
  (* KEEP="TRUE" *) wire n2969_o;
  (* KEEP="TRUE" *) wire n2970_o;
  (* KEEP="TRUE" *) wire n2971_o;
  (* KEEP="TRUE" *) wire n2972_o;
  (* KEEP="TRUE" *) wire n2973_o;
  (* KEEP="TRUE" *) wire n2974_o;
  (* KEEP="TRUE" *) wire n2975_o;
  (* KEEP="TRUE" *) wire n2976_o;
  (* KEEP="TRUE" *) wire n2977_o;
  (* KEEP="TRUE" *) wire n2978_o;
  (* KEEP="TRUE" *) wire n2979_o;
  (* KEEP="TRUE" *) wire n2980_o;
  (* KEEP="TRUE" *) wire n2981_o;
  (* KEEP="TRUE" *) wire n2982_o;
  (* KEEP="TRUE" *) wire n2983_o;
  (* KEEP="TRUE" *) wire n2984_o;
  (* KEEP="TRUE" *) wire n2985_o;
  (* KEEP="TRUE" *) wire n2986_o;
  (* KEEP="TRUE" *) wire n2987_o;
  (* KEEP="TRUE" *) wire n2988_o;
  (* KEEP="TRUE" *) wire n2989_o;
  (* KEEP="TRUE" *) wire n2990_o;
  (* KEEP="TRUE" *) wire n2991_o;
  (* KEEP="TRUE" *) wire n2992_o;
  (* KEEP="TRUE" *) wire n2993_o;
  (* KEEP="TRUE" *) wire n2994_o;
  (* KEEP="TRUE" *) wire n2995_o;
  (* KEEP="TRUE" *) wire n2996_o;
  (* KEEP="TRUE" *) wire n2997_o;
  (* KEEP="TRUE" *) wire n2998_o;
  (* KEEP="TRUE" *) wire n2999_o;
  (* KEEP="TRUE" *) wire n3000_o;
  (* KEEP="TRUE" *) wire n3001_o;
  (* KEEP="TRUE" *) wire n3002_o;
  (* KEEP="TRUE" *) wire n3003_o;
  (* KEEP="TRUE" *) wire n3004_o;
  (* KEEP="TRUE" *) wire n3005_o;
  (* KEEP="TRUE" *) wire n3006_o;
  (* KEEP="TRUE" *) wire n3007_o;
  (* KEEP="TRUE" *) wire n3008_o;
  (* KEEP="TRUE" *) wire n3009_o;
  (* KEEP="TRUE" *) wire n3010_o;
  (* KEEP="TRUE" *) wire n3011_o;
  (* KEEP="TRUE" *) wire n3012_o;
  (* KEEP="TRUE" *) wire n3013_o;
  (* KEEP="TRUE" *) wire n3014_o;
  (* KEEP="TRUE" *) wire n3015_o;
  (* KEEP="TRUE" *) wire n3016_o;
  (* KEEP="TRUE" *) wire n3017_o;
  (* KEEP="TRUE" *) wire n3018_o;
  (* KEEP="TRUE" *) wire n3019_o;
  (* KEEP="TRUE" *) wire n3020_o;
  (* KEEP="TRUE" *) wire n3021_o;
  (* KEEP="TRUE" *) wire n3022_o;
  (* KEEP="TRUE" *) wire n3023_o;
  (* KEEP="TRUE" *) wire n3024_o;
  (* KEEP="TRUE" *) wire n3025_o;
  (* KEEP="TRUE" *) wire n3026_o;
  (* KEEP="TRUE" *) wire n3027_o;
  (* KEEP="TRUE" *) wire n3028_o;
  (* KEEP="TRUE" *) wire n3029_o;
  (* KEEP="TRUE" *) wire n3030_o;
  (* KEEP="TRUE" *) wire n3031_o;
  (* KEEP="TRUE" *) wire n3032_o;
  (* KEEP="TRUE" *) wire n3033_o;
  (* KEEP="TRUE" *) wire n3034_o;
  (* KEEP="TRUE" *) wire n3035_o;
  (* KEEP="TRUE" *) wire n3036_o;
  (* KEEP="TRUE" *) wire n3037_o;
  (* KEEP="TRUE" *) wire n3038_o;
  (* KEEP="TRUE" *) wire n3039_o;
  (* KEEP="TRUE" *) wire n3040_o;
  (* KEEP="TRUE" *) wire n3041_o;
  (* KEEP="TRUE" *) wire n3042_o;
  (* KEEP="TRUE" *) wire n3043_o;
  (* KEEP="TRUE" *) wire n3044_o;
  (* KEEP="TRUE" *) wire n3045_o;
  (* KEEP="TRUE" *) wire n3046_o;
  (* KEEP="TRUE" *) wire n3047_o;
  (* KEEP="TRUE" *) wire n3048_o;
  (* KEEP="TRUE" *) wire n3049_o;
  (* KEEP="TRUE" *) wire n3050_o;
  (* KEEP="TRUE" *) wire n3051_o;
  (* KEEP="TRUE" *) wire n3052_o;
  (* KEEP="TRUE" *) wire n3053_o;
  (* KEEP="TRUE" *) wire n3054_o;
  (* KEEP="TRUE" *) wire n3055_o;
  (* KEEP="TRUE" *) wire n3056_o;
  (* KEEP="TRUE" *) wire n3057_o;
  (* KEEP="TRUE" *) wire n3058_o;
  (* KEEP="TRUE" *) wire n3059_o;
  (* KEEP="TRUE" *) wire n3060_o;
  (* KEEP="TRUE" *) wire n3061_o;
  (* KEEP="TRUE" *) wire n3062_o;
  (* KEEP="TRUE" *) wire n3063_o;
  (* KEEP="TRUE" *) wire n3064_o;
  (* KEEP="TRUE" *) wire n3065_o;
  (* KEEP="TRUE" *) wire n3066_o;
  (* KEEP="TRUE" *) wire n3067_o;
  (* KEEP="TRUE" *) wire n3068_o;
  (* KEEP="TRUE" *) wire n3069_o;
  (* KEEP="TRUE" *) wire n3070_o;
  (* KEEP="TRUE" *) wire n3071_o;
  (* KEEP="TRUE" *) wire n3072_o;
  (* KEEP="TRUE" *) wire n3073_o;
  (* KEEP="TRUE" *) wire n3074_o;
  (* KEEP="TRUE" *) wire n3075_o;
  (* KEEP="TRUE" *) wire n3076_o;
  (* KEEP="TRUE" *) wire n3077_o;
  (* KEEP="TRUE" *) wire n3078_o;
  (* KEEP="TRUE" *) wire n3079_o;
  (* KEEP="TRUE" *) wire n3080_o;
  (* KEEP="TRUE" *) wire n3081_o;
  (* KEEP="TRUE" *) wire n3082_o;
  (* KEEP="TRUE" *) wire n3083_o;
  (* KEEP="TRUE" *) wire n3084_o;
  (* KEEP="TRUE" *) wire n3085_o;
  (* KEEP="TRUE" *) wire n3086_o;
  (* KEEP="TRUE" *) wire n3087_o;
  (* KEEP="TRUE" *) wire n3088_o;
  (* KEEP="TRUE" *) wire n3089_o;
  (* KEEP="TRUE" *) wire n3090_o;
  (* KEEP="TRUE" *) wire n3091_o;
  (* KEEP="TRUE" *) wire n3092_o;
  (* KEEP="TRUE" *) wire n3093_o;
  (* KEEP="TRUE" *) wire n3094_o;
  (* KEEP="TRUE" *) wire n3095_o;
  (* KEEP="TRUE" *) wire n3096_o;
  (* KEEP="TRUE" *) wire n3097_o;
  (* KEEP="TRUE" *) wire n3098_o;
  (* KEEP="TRUE" *) wire n3099_o;
  (* KEEP="TRUE" *) wire n3100_o;
  (* KEEP="TRUE" *) wire n3101_o;
  (* KEEP="TRUE" *) wire n3102_o;
  (* KEEP="TRUE" *) wire n3103_o;
  (* KEEP="TRUE" *) wire n3104_o;
  (* KEEP="TRUE" *) wire n3105_o;
  (* KEEP="TRUE" *) wire n3106_o;
  (* KEEP="TRUE" *) wire n3107_o;
  (* KEEP="TRUE" *) wire n3108_o;
  (* KEEP="TRUE" *) wire n3109_o;
  (* KEEP="TRUE" *) wire n3110_o;
  (* KEEP="TRUE" *) wire n3111_o;
  (* KEEP="TRUE" *) wire n3112_o;
  (* KEEP="TRUE" *) wire n3113_o;
  (* KEEP="TRUE" *) wire n3114_o;
  (* KEEP="TRUE" *) wire n3115_o;
  (* KEEP="TRUE" *) wire n3116_o;
  (* KEEP="TRUE" *) wire n3117_o;
  (* KEEP="TRUE" *) wire n3118_o;
  (* KEEP="TRUE" *) wire n3119_o;
  (* KEEP="TRUE" *) wire n3120_o;
  (* KEEP="TRUE" *) wire n3121_o;
  (* KEEP="TRUE" *) wire n3122_o;
  (* KEEP="TRUE" *) wire n3123_o;
  (* KEEP="TRUE" *) wire n3124_o;
  (* KEEP="TRUE" *) wire n3125_o;
  (* KEEP="TRUE" *) wire n3126_o;
  (* KEEP="TRUE" *) wire n3127_o;
  (* KEEP="TRUE" *) wire n3128_o;
  (* KEEP="TRUE" *) wire n3129_o;
  (* KEEP="TRUE" *) wire n3130_o;
  (* KEEP="TRUE" *) wire n3131_o;
  (* KEEP="TRUE" *) wire n3132_o;
  (* KEEP="TRUE" *) wire n3133_o;
  (* KEEP="TRUE" *) wire n3134_o;
  (* KEEP="TRUE" *) wire n3135_o;
  (* KEEP="TRUE" *) wire n3136_o;
  (* KEEP="TRUE" *) wire n3137_o;
  (* KEEP="TRUE" *) wire n3138_o;
  (* KEEP="TRUE" *) wire n3139_o;
  (* KEEP="TRUE" *) wire n3140_o;
  (* KEEP="TRUE" *) wire n3141_o;
  (* KEEP="TRUE" *) wire n3142_o;
  (* KEEP="TRUE" *) wire n3143_o;
  (* KEEP="TRUE" *) wire n3144_o;
  (* KEEP="TRUE" *) wire n3145_o;
  (* KEEP="TRUE" *) wire n3146_o;
  (* KEEP="TRUE" *) wire n3147_o;
  (* KEEP="TRUE" *) wire n3148_o;
  (* KEEP="TRUE" *) wire n3149_o;
  (* KEEP="TRUE" *) wire n3150_o;
  (* KEEP="TRUE" *) wire n3151_o;
  (* KEEP="TRUE" *) wire n3152_o;
  (* KEEP="TRUE" *) wire n3153_o;
  (* KEEP="TRUE" *) wire n3154_o;
  (* KEEP="TRUE" *) wire n3155_o;
  (* KEEP="TRUE" *) wire n3156_o;
  (* KEEP="TRUE" *) wire n3157_o;
  (* KEEP="TRUE" *) wire n3158_o;
  (* KEEP="TRUE" *) wire n3159_o;
  (* KEEP="TRUE" *) wire n3160_o;
  (* KEEP="TRUE" *) wire n3161_o;
  (* KEEP="TRUE" *) wire n3162_o;
  (* KEEP="TRUE" *) wire n3163_o;
  (* KEEP="TRUE" *) wire n3164_o;
  (* KEEP="TRUE" *) wire n3165_o;
  (* KEEP="TRUE" *) wire n3166_o;
  (* KEEP="TRUE" *) wire n3167_o;
  (* KEEP="TRUE" *) wire n3168_o;
  (* KEEP="TRUE" *) wire n3169_o;
  (* KEEP="TRUE" *) wire n3170_o;
  (* KEEP="TRUE" *) wire n3171_o;
  (* KEEP="TRUE" *) wire n3172_o;
  (* KEEP="TRUE" *) wire n3173_o;
  (* KEEP="TRUE" *) wire n3174_o;
  (* KEEP="TRUE" *) wire n3175_o;
  (* KEEP="TRUE" *) wire n3176_o;
  (* KEEP="TRUE" *) wire n3177_o;
  (* KEEP="TRUE" *) wire n3178_o;
  (* KEEP="TRUE" *) wire n3179_o;
  (* KEEP="TRUE" *) wire n3180_o;
  (* KEEP="TRUE" *) wire n3181_o;
  (* KEEP="TRUE" *) wire n3182_o;
  (* KEEP="TRUE" *) wire n3183_o;
  (* KEEP="TRUE" *) wire n3184_o;
  (* KEEP="TRUE" *) wire n3185_o;
  (* KEEP="TRUE" *) wire n3186_o;
  (* KEEP="TRUE" *) wire n3187_o;
  (* KEEP="TRUE" *) wire n3188_o;
  (* KEEP="TRUE" *) wire n3189_o;
  (* KEEP="TRUE" *) wire n3190_o;
  (* KEEP="TRUE" *) wire n3191_o;
  (* KEEP="TRUE" *) wire n3192_o;
  (* KEEP="TRUE" *) wire n3193_o;
  (* KEEP="TRUE" *) wire n3194_o;
  (* KEEP="TRUE" *) wire n3195_o;
  (* KEEP="TRUE" *) wire n3196_o;
  (* KEEP="TRUE" *) wire n3197_o;
  (* KEEP="TRUE" *) wire n3198_o;
  (* KEEP="TRUE" *) wire n3199_o;
  (* KEEP="TRUE" *) wire n3200_o;
  (* KEEP="TRUE" *) wire n3201_o;
  (* KEEP="TRUE" *) wire n3202_o;
  (* KEEP="TRUE" *) wire n3203_o;
  (* KEEP="TRUE" *) wire n3204_o;
  (* KEEP="TRUE" *) wire n3205_o;
  (* KEEP="TRUE" *) wire n3206_o;
  (* KEEP="TRUE" *) wire n3207_o;
  (* KEEP="TRUE" *) wire n3208_o;
  (* KEEP="TRUE" *) wire n3209_o;
  (* KEEP="TRUE" *) wire n3210_o;
  (* KEEP="TRUE" *) wire n3211_o;
  (* KEEP="TRUE" *) wire n3212_o;
  (* KEEP="TRUE" *) wire n3213_o;
  (* KEEP="TRUE" *) wire n3214_o;
  (* KEEP="TRUE" *) wire n3215_o;
  (* KEEP="TRUE" *) wire n3216_o;
  (* KEEP="TRUE" *) wire n3217_o;
  (* KEEP="TRUE" *) wire n3218_o;
  (* KEEP="TRUE" *) wire n3219_o;
  (* KEEP="TRUE" *) wire n3220_o;
  (* KEEP="TRUE" *) wire n3221_o;
  (* KEEP="TRUE" *) wire n3222_o;
  (* KEEP="TRUE" *) wire n3223_o;
  (* KEEP="TRUE" *) wire n3224_o;
  (* KEEP="TRUE" *) wire n3225_o;
  (* KEEP="TRUE" *) wire n3226_o;
  (* KEEP="TRUE" *) wire n3227_o;
  (* KEEP="TRUE" *) wire n3228_o;
  (* KEEP="TRUE" *) wire n3229_o;
  (* KEEP="TRUE" *) wire n3230_o;
  (* KEEP="TRUE" *) wire n3231_o;
  (* KEEP="TRUE" *) wire n3232_o;
  (* KEEP="TRUE" *) wire n3233_o;
  (* KEEP="TRUE" *) wire n3234_o;
  (* KEEP="TRUE" *) wire n3235_o;
  (* KEEP="TRUE" *) wire n3236_o;
  (* KEEP="TRUE" *) wire n3237_o;
  (* KEEP="TRUE" *) wire n3238_o;
  (* KEEP="TRUE" *) wire n3239_o;
  (* KEEP="TRUE" *) wire n3240_o;
  (* KEEP="TRUE" *) wire n3241_o;
  (* KEEP="TRUE" *) wire n3242_o;
  (* KEEP="TRUE" *) wire n3243_o;
  (* KEEP="TRUE" *) wire n3244_o;
  (* KEEP="TRUE" *) wire n3245_o;
  (* KEEP="TRUE" *) wire n3246_o;
  (* KEEP="TRUE" *) wire n3247_o;
  (* KEEP="TRUE" *) wire n3248_o;
  (* KEEP="TRUE" *) wire n3249_o;
  (* KEEP="TRUE" *) wire n3250_o;
  (* KEEP="TRUE" *) wire n3251_o;
  (* KEEP="TRUE" *) wire n3252_o;
  (* KEEP="TRUE" *) wire n3253_o;
  (* KEEP="TRUE" *) wire n3254_o;
  (* KEEP="TRUE" *) wire n3255_o;
  (* KEEP="TRUE" *) wire n3256_o;
  (* KEEP="TRUE" *) wire n3257_o;
  (* KEEP="TRUE" *) wire n3258_o;
  (* KEEP="TRUE" *) wire n3259_o;
  (* KEEP="TRUE" *) wire n3260_o;
  (* KEEP="TRUE" *) wire n3261_o;
  (* KEEP="TRUE" *) wire n3262_o;
  (* KEEP="TRUE" *) wire n3263_o;
  (* KEEP="TRUE" *) wire n3264_o;
  (* KEEP="TRUE" *) wire n3265_o;
  (* KEEP="TRUE" *) wire n3266_o;
  (* KEEP="TRUE" *) wire n3267_o;
  (* KEEP="TRUE" *) wire n3268_o;
  (* KEEP="TRUE" *) wire n3269_o;
  (* KEEP="TRUE" *) wire n3270_o;
  (* KEEP="TRUE" *) wire n3271_o;
  (* KEEP="TRUE" *) wire n3272_o;
  (* KEEP="TRUE" *) wire n3273_o;
  (* KEEP="TRUE" *) wire n3274_o;
  (* KEEP="TRUE" *) wire n3275_o;
  (* KEEP="TRUE" *) wire n3276_o;
  (* KEEP="TRUE" *) wire n3277_o;
  (* KEEP="TRUE" *) wire n3278_o;
  (* KEEP="TRUE" *) wire n3279_o;
  (* KEEP="TRUE" *) wire n3280_o;
  (* KEEP="TRUE" *) wire n3281_o;
  (* KEEP="TRUE" *) wire n3282_o;
  (* KEEP="TRUE" *) wire n3283_o;
  (* KEEP="TRUE" *) wire n3284_o;
  (* KEEP="TRUE" *) wire n3285_o;
  (* KEEP="TRUE" *) wire n3286_o;
  (* KEEP="TRUE" *) wire n3287_o;
  (* KEEP="TRUE" *) wire n3288_o;
  (* KEEP="TRUE" *) wire n3289_o;
  (* KEEP="TRUE" *) wire n3290_o;
  (* KEEP="TRUE" *) wire n3291_o;
  (* KEEP="TRUE" *) wire n3292_o;
  (* KEEP="TRUE" *) wire n3293_o;
  (* KEEP="TRUE" *) wire n3294_o;
  (* KEEP="TRUE" *) wire n3295_o;
  (* KEEP="TRUE" *) wire n3296_o;
  (* KEEP="TRUE" *) wire n3297_o;
  (* KEEP="TRUE" *) wire n3298_o;
  (* KEEP="TRUE" *) wire n3299_o;
  (* KEEP="TRUE" *) wire n3300_o;
  (* KEEP="TRUE" *) wire n3301_o;
  (* KEEP="TRUE" *) wire n3302_o;
  (* KEEP="TRUE" *) wire n3303_o;
  (* KEEP="TRUE" *) wire n3304_o;
  (* KEEP="TRUE" *) wire n3305_o;
  (* KEEP="TRUE" *) wire n3306_o;
  (* KEEP="TRUE" *) wire n3307_o;
  (* KEEP="TRUE" *) wire n3308_o;
  (* KEEP="TRUE" *) wire n3309_o;
  (* KEEP="TRUE" *) wire n3310_o;
  (* KEEP="TRUE" *) wire n3311_o;
  (* KEEP="TRUE" *) wire n3312_o;
  (* KEEP="TRUE" *) wire n3313_o;
  (* KEEP="TRUE" *) wire n3314_o;
  (* KEEP="TRUE" *) wire n3315_o;
  (* KEEP="TRUE" *) wire n3316_o;
  (* KEEP="TRUE" *) wire n3317_o;
  (* KEEP="TRUE" *) wire n3318_o;
  (* KEEP="TRUE" *) wire n3319_o;
  (* KEEP="TRUE" *) wire n3320_o;
  (* KEEP="TRUE" *) wire n3321_o;
  (* KEEP="TRUE" *) wire n3322_o;
  (* KEEP="TRUE" *) wire n3323_o;
  (* KEEP="TRUE" *) wire n3324_o;
  (* KEEP="TRUE" *) wire n3325_o;
  (* KEEP="TRUE" *) wire n3326_o;
  (* KEEP="TRUE" *) wire n3327_o;
  (* KEEP="TRUE" *) wire n3328_o;
  (* KEEP="TRUE" *) wire n3329_o;
  (* KEEP="TRUE" *) wire n3330_o;
  (* KEEP="TRUE" *) wire n3331_o;
  (* KEEP="TRUE" *) wire n3332_o;
  (* KEEP="TRUE" *) wire n3333_o;
  (* KEEP="TRUE" *) wire n3334_o;
  (* KEEP="TRUE" *) wire n3335_o;
  (* KEEP="TRUE" *) wire n3336_o;
  (* KEEP="TRUE" *) wire n3337_o;
  (* KEEP="TRUE" *) wire n3338_o;
  (* KEEP="TRUE" *) wire n3339_o;
  (* KEEP="TRUE" *) wire n3340_o;
  (* KEEP="TRUE" *) wire n3341_o;
  (* KEEP="TRUE" *) wire n3342_o;
  (* KEEP="TRUE" *) wire n3343_o;
  (* KEEP="TRUE" *) wire n3344_o;
  (* KEEP="TRUE" *) wire n3345_o;
  (* KEEP="TRUE" *) wire n3346_o;
  (* KEEP="TRUE" *) wire n3347_o;
  (* KEEP="TRUE" *) wire n3348_o;
  (* KEEP="TRUE" *) wire n3349_o;
  (* KEEP="TRUE" *) wire n3350_o;
  (* KEEP="TRUE" *) wire n3351_o;
  (* KEEP="TRUE" *) wire n3352_o;
  (* KEEP="TRUE" *) wire n3353_o;
  (* KEEP="TRUE" *) wire n3354_o;
  (* KEEP="TRUE" *) wire n3355_o;
  (* KEEP="TRUE" *) wire n3356_o;
  (* KEEP="TRUE" *) wire n3357_o;
  (* KEEP="TRUE" *) wire n3358_o;
  (* KEEP="TRUE" *) wire n3359_o;
  (* KEEP="TRUE" *) wire n3360_o;
  (* KEEP="TRUE" *) wire n3361_o;
  (* KEEP="TRUE" *) wire n3362_o;
  (* KEEP="TRUE" *) wire n3363_o;
  (* KEEP="TRUE" *) wire n3364_o;
  (* KEEP="TRUE" *) wire n3365_o;
  (* KEEP="TRUE" *) wire n3366_o;
  (* KEEP="TRUE" *) wire n3367_o;
  (* KEEP="TRUE" *) wire n3368_o;
  (* KEEP="TRUE" *) wire n3369_o;
  (* KEEP="TRUE" *) wire n3370_o;
  (* KEEP="TRUE" *) wire n3371_o;
  (* KEEP="TRUE" *) wire n3372_o;
  (* KEEP="TRUE" *) wire n3373_o;
  (* KEEP="TRUE" *) wire n3374_o;
  (* KEEP="TRUE" *) wire n3375_o;
  (* KEEP="TRUE" *) wire n3376_o;
  (* KEEP="TRUE" *) wire n3377_o;
  (* KEEP="TRUE" *) wire n3378_o;
  (* KEEP="TRUE" *) wire n3379_o;
  (* KEEP="TRUE" *) wire n3380_o;
  (* KEEP="TRUE" *) wire n3381_o;
  (* KEEP="TRUE" *) wire n3382_o;
  (* KEEP="TRUE" *) wire n3383_o;
  (* KEEP="TRUE" *) wire n3384_o;
  (* KEEP="TRUE" *) wire n3385_o;
  (* KEEP="TRUE" *) wire n3386_o;
  (* KEEP="TRUE" *) wire n3387_o;
  (* KEEP="TRUE" *) wire n3388_o;
  (* KEEP="TRUE" *) wire n3389_o;
  (* KEEP="TRUE" *) wire n3390_o;
  (* KEEP="TRUE" *) wire n3391_o;
  (* KEEP="TRUE" *) wire n3392_o;
  (* KEEP="TRUE" *) wire n3393_o;
  (* KEEP="TRUE" *) wire n3394_o;
  (* KEEP="TRUE" *) wire n3395_o;
  (* KEEP="TRUE" *) wire n3396_o;
  (* KEEP="TRUE" *) wire n3397_o;
  (* KEEP="TRUE" *) wire n3398_o;
  (* KEEP="TRUE" *) wire n3399_o;
  (* KEEP="TRUE" *) wire n3400_o;
  (* KEEP="TRUE" *) wire n3401_o;
  (* KEEP="TRUE" *) wire n3402_o;
  (* KEEP="TRUE" *) wire n3403_o;
  (* KEEP="TRUE" *) wire n3404_o;
  (* KEEP="TRUE" *) wire n3405_o;
  (* KEEP="TRUE" *) wire n3406_o;
  (* KEEP="TRUE" *) wire n3407_o;
  (* KEEP="TRUE" *) wire n3408_o;
  (* KEEP="TRUE" *) wire n3409_o;
  (* KEEP="TRUE" *) wire n3410_o;
  (* KEEP="TRUE" *) wire n3411_o;
  (* KEEP="TRUE" *) wire n3412_o;
  (* KEEP="TRUE" *) wire n3413_o;
  (* KEEP="TRUE" *) wire n3414_o;
  (* KEEP="TRUE" *) wire n3415_o;
  (* KEEP="TRUE" *) wire n3416_o;
  (* KEEP="TRUE" *) wire n3417_o;
  (* KEEP="TRUE" *) wire n3418_o;
  (* KEEP="TRUE" *) wire n3419_o;
  (* KEEP="TRUE" *) wire n3420_o;
  (* KEEP="TRUE" *) wire n3421_o;
  (* KEEP="TRUE" *) wire n3422_o;
  (* KEEP="TRUE" *) wire n3423_o;
  (* KEEP="TRUE" *) wire n3424_o;
  (* KEEP="TRUE" *) wire n3425_o;
  (* KEEP="TRUE" *) wire n3426_o;
  (* KEEP="TRUE" *) wire n3427_o;
  (* KEEP="TRUE" *) wire n3428_o;
  (* KEEP="TRUE" *) wire n3429_o;
  (* KEEP="TRUE" *) wire n3430_o;
  (* KEEP="TRUE" *) wire n3431_o;
  (* KEEP="TRUE" *) wire n3432_o;
  (* KEEP="TRUE" *) wire n3433_o;
  (* KEEP="TRUE" *) wire n3434_o;
  (* KEEP="TRUE" *) wire n3435_o;
  (* KEEP="TRUE" *) wire n3436_o;
  (* KEEP="TRUE" *) wire n3437_o;
  (* KEEP="TRUE" *) wire n3438_o;
  (* KEEP="TRUE" *) wire n3439_o;
  (* KEEP="TRUE" *) wire n3440_o;
  (* KEEP="TRUE" *) wire n3441_o;
  (* KEEP="TRUE" *) wire n3442_o;
  (* KEEP="TRUE" *) wire n3443_o;
  (* KEEP="TRUE" *) wire n3444_o;
  (* KEEP="TRUE" *) wire n3445_o;
  (* KEEP="TRUE" *) wire n3446_o;
  (* KEEP="TRUE" *) wire n3447_o;
  (* KEEP="TRUE" *) wire n3448_o;
  (* KEEP="TRUE" *) wire n3449_o;
  (* KEEP="TRUE" *) wire n3450_o;
  (* KEEP="TRUE" *) wire n3451_o;
  (* KEEP="TRUE" *) wire n3452_o;
  (* KEEP="TRUE" *) wire n3453_o;
  (* KEEP="TRUE" *) wire n3454_o;
  (* KEEP="TRUE" *) wire n3455_o;
  (* KEEP="TRUE" *) wire n3456_o;
  (* KEEP="TRUE" *) wire n3457_o;
  (* KEEP="TRUE" *) wire n3458_o;
  (* KEEP="TRUE" *) wire n3459_o;
  (* KEEP="TRUE" *) wire n3460_o;
  (* KEEP="TRUE" *) wire n3461_o;
  (* KEEP="TRUE" *) wire n3462_o;
  (* KEEP="TRUE" *) wire n3463_o;
  (* KEEP="TRUE" *) wire n3464_o;
  (* KEEP="TRUE" *) wire n3465_o;
  (* KEEP="TRUE" *) wire n3466_o;
  (* KEEP="TRUE" *) wire n3467_o;
  (* KEEP="TRUE" *) wire n3468_o;
  (* KEEP="TRUE" *) wire n3469_o;
  (* KEEP="TRUE" *) wire n3470_o;
  (* KEEP="TRUE" *) wire n3471_o;
  (* KEEP="TRUE" *) wire n3472_o;
  (* KEEP="TRUE" *) wire n3473_o;
  (* KEEP="TRUE" *) wire n3474_o;
  (* KEEP="TRUE" *) wire n3475_o;
  (* KEEP="TRUE" *) wire n3476_o;
  (* KEEP="TRUE" *) wire n3477_o;
  (* KEEP="TRUE" *) wire n3478_o;
  (* KEEP="TRUE" *) wire n3479_o;
  (* KEEP="TRUE" *) wire n3480_o;
  (* KEEP="TRUE" *) wire n3481_o;
  (* KEEP="TRUE" *) wire n3482_o;
  (* KEEP="TRUE" *) wire n3483_o;
  (* KEEP="TRUE" *) wire n3484_o;
  (* KEEP="TRUE" *) wire n3485_o;
  (* KEEP="TRUE" *) wire n3486_o;
  (* KEEP="TRUE" *) wire n3487_o;
  (* KEEP="TRUE" *) wire n3488_o;
  (* KEEP="TRUE" *) wire n3489_o;
  (* KEEP="TRUE" *) wire n3490_o;
  (* KEEP="TRUE" *) wire n3491_o;
  (* KEEP="TRUE" *) wire n3492_o;
  (* KEEP="TRUE" *) wire n3493_o;
  (* KEEP="TRUE" *) wire n3494_o;
  (* KEEP="TRUE" *) wire n3495_o;
  (* KEEP="TRUE" *) wire n3496_o;
  (* KEEP="TRUE" *) wire n3497_o;
  (* KEEP="TRUE" *) wire n3498_o;
  (* KEEP="TRUE" *) wire n3499_o;
  (* KEEP="TRUE" *) wire n3500_o;
  (* KEEP="TRUE" *) wire n3501_o;
  (* KEEP="TRUE" *) wire n3502_o;
  (* KEEP="TRUE" *) wire n3503_o;
  (* KEEP="TRUE" *) wire n3504_o;
  (* KEEP="TRUE" *) wire n3505_o;
  (* KEEP="TRUE" *) wire n3506_o;
  (* KEEP="TRUE" *) wire n3507_o;
  (* KEEP="TRUE" *) wire n3508_o;
  (* KEEP="TRUE" *) wire n3509_o;
  (* KEEP="TRUE" *) wire n3510_o;
  (* KEEP="TRUE" *) wire n3511_o;
  (* KEEP="TRUE" *) wire n3512_o;
  (* KEEP="TRUE" *) wire n3513_o;
  (* KEEP="TRUE" *) wire n3514_o;
  (* KEEP="TRUE" *) wire n3515_o;
  (* KEEP="TRUE" *) wire n3516_o;
  (* KEEP="TRUE" *) wire n3517_o;
  (* KEEP="TRUE" *) wire n3518_o;
  (* KEEP="TRUE" *) wire n3519_o;
  (* KEEP="TRUE" *) wire n3520_o;
  (* KEEP="TRUE" *) wire n3521_o;
  (* KEEP="TRUE" *) wire n3522_o;
  (* KEEP="TRUE" *) wire n3523_o;
  (* KEEP="TRUE" *) wire n3524_o;
  (* KEEP="TRUE" *) wire n3525_o;
  (* KEEP="TRUE" *) wire n3526_o;
  (* KEEP="TRUE" *) wire n3527_o;
  (* KEEP="TRUE" *) wire n3528_o;
  (* KEEP="TRUE" *) wire n3529_o;
  (* KEEP="TRUE" *) wire n3530_o;
  (* KEEP="TRUE" *) wire n3531_o;
  (* KEEP="TRUE" *) wire n3532_o;
  (* KEEP="TRUE" *) wire n3533_o;
  (* KEEP="TRUE" *) wire n3534_o;
  (* KEEP="TRUE" *) wire n3535_o;
  (* KEEP="TRUE" *) wire n3536_o;
  (* KEEP="TRUE" *) wire n3537_o;
  (* KEEP="TRUE" *) wire n3538_o;
  (* KEEP="TRUE" *) wire n3539_o;
  (* KEEP="TRUE" *) wire n3540_o;
  (* KEEP="TRUE" *) wire n3541_o;
  (* KEEP="TRUE" *) wire n3542_o;
  (* KEEP="TRUE" *) wire n3543_o;
  (* KEEP="TRUE" *) wire n3544_o;
  (* KEEP="TRUE" *) wire n3545_o;
  (* KEEP="TRUE" *) wire n3546_o;
  (* KEEP="TRUE" *) wire n3547_o;
  (* KEEP="TRUE" *) wire n3548_o;
  (* KEEP="TRUE" *) wire n3549_o;
  (* KEEP="TRUE" *) wire n3550_o;
  (* KEEP="TRUE" *) wire n3551_o;
  (* KEEP="TRUE" *) wire n3552_o;
  (* KEEP="TRUE" *) wire n3553_o;
  (* KEEP="TRUE" *) wire n3554_o;
  (* KEEP="TRUE" *) wire n3555_o;
  (* KEEP="TRUE" *) wire n3556_o;
  (* KEEP="TRUE" *) wire n3557_o;
  (* KEEP="TRUE" *) wire n3558_o;
  (* KEEP="TRUE" *) wire n3559_o;
  (* KEEP="TRUE" *) wire n3560_o;
  (* KEEP="TRUE" *) wire n3561_o;
  (* KEEP="TRUE" *) wire n3562_o;
  (* KEEP="TRUE" *) wire n3563_o;
  (* KEEP="TRUE" *) wire n3564_o;
  (* KEEP="TRUE" *) wire n3565_o;
  (* KEEP="TRUE" *) wire n3566_o;
  (* KEEP="TRUE" *) wire n3567_o;
  (* KEEP="TRUE" *) wire n3568_o;
  (* KEEP="TRUE" *) wire n3569_o;
  (* KEEP="TRUE" *) wire n3570_o;
  (* KEEP="TRUE" *) wire n3571_o;
  (* KEEP="TRUE" *) wire n3572_o;
  (* KEEP="TRUE" *) wire n3573_o;
  (* KEEP="TRUE" *) wire n3574_o;
  (* KEEP="TRUE" *) wire n3575_o;
  (* KEEP="TRUE" *) wire n3576_o;
  (* KEEP="TRUE" *) wire n3577_o;
  (* KEEP="TRUE" *) wire n3578_o;
  (* KEEP="TRUE" *) wire n3579_o;
  (* KEEP="TRUE" *) wire n3580_o;
  (* KEEP="TRUE" *) wire n3581_o;
  (* KEEP="TRUE" *) wire n3582_o;
  (* KEEP="TRUE" *) wire n3583_o;
  (* KEEP="TRUE" *) wire n3584_o;
  (* KEEP="TRUE" *) wire n3585_o;
  (* KEEP="TRUE" *) wire n3586_o;
  (* KEEP="TRUE" *) wire n3587_o;
  (* KEEP="TRUE" *) wire n3588_o;
  (* KEEP="TRUE" *) wire n3589_o;
  (* KEEP="TRUE" *) wire n3590_o;
  (* KEEP="TRUE" *) wire n3591_o;
  (* KEEP="TRUE" *) wire n3592_o;
  (* KEEP="TRUE" *) wire n3593_o;
  (* KEEP="TRUE" *) wire n3594_o;
  (* KEEP="TRUE" *) wire n3595_o;
  (* KEEP="TRUE" *) wire n3596_o;
  (* KEEP="TRUE" *) wire n3597_o;
  (* KEEP="TRUE" *) wire n3598_o;
  (* KEEP="TRUE" *) wire n3599_o;
  (* KEEP="TRUE" *) wire n3600_o;
  (* KEEP="TRUE" *) wire n3601_o;
  (* KEEP="TRUE" *) wire n3602_o;
  (* KEEP="TRUE" *) wire n3603_o;
  (* KEEP="TRUE" *) wire n3604_o;
  (* KEEP="TRUE" *) wire n3605_o;
  (* KEEP="TRUE" *) wire n3606_o;
  (* KEEP="TRUE" *) wire [255:0] n3607_o;
  (* KEEP="TRUE" *) wire n3608_o;
  (* KEEP="TRUE" *) wire n3609_o;
  (* KEEP="TRUE" *) wire n3610_o;
  (* KEEP="TRUE" *) wire n3611_o;
  (* KEEP="TRUE" *) wire n3612_o;
  (* KEEP="TRUE" *) wire n3613_o;
  (* KEEP="TRUE" *) wire n3614_o;
  (* KEEP="TRUE" *) wire n3615_o;
  (* KEEP="TRUE" *) wire n3616_o;
  (* KEEP="TRUE" *) wire n3617_o;
  (* KEEP="TRUE" *) wire n3618_o;
  (* KEEP="TRUE" *) wire n3619_o;
  (* KEEP="TRUE" *) wire n3620_o;
  (* KEEP="TRUE" *) wire n3621_o;
  (* KEEP="TRUE" *) wire n3622_o;
  (* KEEP="TRUE" *) wire n3623_o;
  (* KEEP="TRUE" *) wire n3624_o;
  (* KEEP="TRUE" *) wire n3625_o;
  (* KEEP="TRUE" *) wire n3626_o;
  (* KEEP="TRUE" *) wire n3627_o;
  (* KEEP="TRUE" *) wire n3628_o;
  (* KEEP="TRUE" *) wire n3629_o;
  (* KEEP="TRUE" *) wire n3630_o;
  (* KEEP="TRUE" *) wire n3631_o;
  (* KEEP="TRUE" *) wire n3632_o;
  (* KEEP="TRUE" *) wire n3633_o;
  (* KEEP="TRUE" *) wire n3634_o;
  (* KEEP="TRUE" *) wire n3635_o;
  (* KEEP="TRUE" *) wire n3636_o;
  (* KEEP="TRUE" *) wire n3637_o;
  (* KEEP="TRUE" *) wire n3638_o;
  (* KEEP="TRUE" *) wire n3639_o;
  (* KEEP="TRUE" *) wire n3640_o;
  (* KEEP="TRUE" *) wire n3641_o;
  (* KEEP="TRUE" *) wire n3642_o;
  (* KEEP="TRUE" *) wire n3643_o;
  (* KEEP="TRUE" *) wire n3644_o;
  (* KEEP="TRUE" *) wire n3645_o;
  (* KEEP="TRUE" *) wire n3646_o;
  (* KEEP="TRUE" *) wire n3647_o;
  (* KEEP="TRUE" *) wire n3648_o;
  (* KEEP="TRUE" *) wire n3649_o;
  (* KEEP="TRUE" *) wire n3650_o;
  (* KEEP="TRUE" *) wire n3651_o;
  (* KEEP="TRUE" *) wire n3652_o;
  (* KEEP="TRUE" *) wire n3653_o;
  (* KEEP="TRUE" *) wire n3654_o;
  (* KEEP="TRUE" *) wire n3655_o;
  (* KEEP="TRUE" *) wire n3656_o;
  (* KEEP="TRUE" *) wire n3657_o;
  (* KEEP="TRUE" *) wire n3658_o;
  (* KEEP="TRUE" *) wire n3659_o;
  (* KEEP="TRUE" *) wire n3660_o;
  (* KEEP="TRUE" *) wire n3661_o;
  (* KEEP="TRUE" *) wire n3662_o;
  (* KEEP="TRUE" *) wire n3663_o;
  (* KEEP="TRUE" *) wire n3664_o;
  (* KEEP="TRUE" *) wire n3665_o;
  (* KEEP="TRUE" *) wire n3666_o;
  (* KEEP="TRUE" *) wire n3667_o;
  (* KEEP="TRUE" *) wire n3668_o;
  (* KEEP="TRUE" *) wire n3669_o;
  (* KEEP="TRUE" *) wire n3670_o;
  (* KEEP="TRUE" *) wire n3671_o;
  (* KEEP="TRUE" *) wire n3672_o;
  (* KEEP="TRUE" *) wire n3673_o;
  (* KEEP="TRUE" *) wire n3674_o;
  (* KEEP="TRUE" *) wire n3675_o;
  (* KEEP="TRUE" *) wire n3676_o;
  (* KEEP="TRUE" *) wire n3677_o;
  (* KEEP="TRUE" *) wire n3678_o;
  (* KEEP="TRUE" *) wire n3679_o;
  (* KEEP="TRUE" *) wire n3680_o;
  (* KEEP="TRUE" *) wire n3681_o;
  (* KEEP="TRUE" *) wire n3682_o;
  (* KEEP="TRUE" *) wire n3683_o;
  (* KEEP="TRUE" *) wire n3684_o;
  (* KEEP="TRUE" *) wire n3685_o;
  (* KEEP="TRUE" *) wire n3686_o;
  (* KEEP="TRUE" *) wire n3687_o;
  (* KEEP="TRUE" *) wire n3688_o;
  (* KEEP="TRUE" *) wire n3689_o;
  (* KEEP="TRUE" *) wire n3690_o;
  (* KEEP="TRUE" *) wire n3691_o;
  (* KEEP="TRUE" *) wire n3692_o;
  (* KEEP="TRUE" *) wire n3693_o;
  (* KEEP="TRUE" *) wire n3694_o;
  (* KEEP="TRUE" *) wire n3695_o;
  (* KEEP="TRUE" *) wire n3696_o;
  (* KEEP="TRUE" *) wire n3697_o;
  (* KEEP="TRUE" *) wire n3698_o;
  (* KEEP="TRUE" *) wire n3699_o;
  (* KEEP="TRUE" *) wire n3700_o;
  (* KEEP="TRUE" *) wire n3701_o;
  (* KEEP="TRUE" *) wire n3702_o;
  (* KEEP="TRUE" *) wire n3703_o;
  (* KEEP="TRUE" *) wire n3704_o;
  (* KEEP="TRUE" *) wire n3705_o;
  (* KEEP="TRUE" *) wire n3706_o;
  (* KEEP="TRUE" *) wire n3707_o;
  (* KEEP="TRUE" *) wire n3708_o;
  (* KEEP="TRUE" *) wire n3709_o;
  (* KEEP="TRUE" *) wire n3710_o;
  (* KEEP="TRUE" *) wire n3711_o;
  (* KEEP="TRUE" *) wire n3712_o;
  (* KEEP="TRUE" *) wire n3713_o;
  (* KEEP="TRUE" *) wire n3714_o;
  (* KEEP="TRUE" *) wire n3715_o;
  (* KEEP="TRUE" *) wire n3716_o;
  (* KEEP="TRUE" *) wire n3717_o;
  (* KEEP="TRUE" *) wire n3718_o;
  (* KEEP="TRUE" *) wire n3719_o;
  (* KEEP="TRUE" *) wire n3720_o;
  (* KEEP="TRUE" *) wire n3721_o;
  (* KEEP="TRUE" *) wire n3722_o;
  (* KEEP="TRUE" *) wire n3723_o;
  (* KEEP="TRUE" *) wire n3724_o;
  (* KEEP="TRUE" *) wire n3725_o;
  (* KEEP="TRUE" *) wire n3726_o;
  (* KEEP="TRUE" *) wire n3727_o;
  (* KEEP="TRUE" *) wire n3728_o;
  (* KEEP="TRUE" *) wire n3729_o;
  (* KEEP="TRUE" *) wire n3730_o;
  (* KEEP="TRUE" *) wire n3731_o;
  (* KEEP="TRUE" *) wire n3732_o;
  (* KEEP="TRUE" *) wire n3733_o;
  (* KEEP="TRUE" *) wire n3734_o;
  (* KEEP="TRUE" *) wire n3735_o;
  (* KEEP="TRUE" *) wire n3736_o;
  (* KEEP="TRUE" *) wire n3737_o;
  (* KEEP="TRUE" *) wire n3738_o;
  (* KEEP="TRUE" *) wire n3739_o;
  (* KEEP="TRUE" *) wire n3740_o;
  (* KEEP="TRUE" *) wire n3741_o;
  (* KEEP="TRUE" *) wire n3742_o;
  (* KEEP="TRUE" *) wire n3743_o;
  (* KEEP="TRUE" *) wire n3744_o;
  (* KEEP="TRUE" *) wire n3745_o;
  (* KEEP="TRUE" *) wire n3746_o;
  (* KEEP="TRUE" *) wire n3747_o;
  (* KEEP="TRUE" *) wire n3748_o;
  (* KEEP="TRUE" *) wire n3749_o;
  (* KEEP="TRUE" *) wire n3750_o;
  (* KEEP="TRUE" *) wire n3751_o;
  (* KEEP="TRUE" *) wire n3752_o;
  (* KEEP="TRUE" *) wire n3753_o;
  (* KEEP="TRUE" *) wire n3754_o;
  (* KEEP="TRUE" *) wire n3755_o;
  (* KEEP="TRUE" *) wire n3756_o;
  (* KEEP="TRUE" *) wire n3757_o;
  (* KEEP="TRUE" *) wire n3758_o;
  (* KEEP="TRUE" *) wire n3759_o;
  (* KEEP="TRUE" *) wire n3760_o;
  (* KEEP="TRUE" *) wire n3761_o;
  (* KEEP="TRUE" *) wire n3762_o;
  (* KEEP="TRUE" *) wire n3763_o;
  (* KEEP="TRUE" *) wire n3764_o;
  (* KEEP="TRUE" *) wire n3765_o;
  (* KEEP="TRUE" *) wire n3766_o;
  (* KEEP="TRUE" *) wire n3767_o;
  (* KEEP="TRUE" *) wire n3768_o;
  (* KEEP="TRUE" *) wire n3769_o;
  (* KEEP="TRUE" *) wire n3770_o;
  (* KEEP="TRUE" *) wire n3771_o;
  (* KEEP="TRUE" *) wire n3772_o;
  (* KEEP="TRUE" *) wire n3773_o;
  (* KEEP="TRUE" *) wire n3774_o;
  (* KEEP="TRUE" *) wire n3775_o;
  (* KEEP="TRUE" *) wire n3776_o;
  (* KEEP="TRUE" *) wire n3777_o;
  (* KEEP="TRUE" *) wire n3778_o;
  (* KEEP="TRUE" *) wire n3779_o;
  (* KEEP="TRUE" *) wire n3780_o;
  (* KEEP="TRUE" *) wire n3781_o;
  (* KEEP="TRUE" *) wire n3782_o;
  (* KEEP="TRUE" *) wire n3783_o;
  (* KEEP="TRUE" *) wire n3784_o;
  (* KEEP="TRUE" *) wire n3785_o;
  (* KEEP="TRUE" *) wire n3786_o;
  (* KEEP="TRUE" *) wire n3787_o;
  (* KEEP="TRUE" *) wire n3788_o;
  (* KEEP="TRUE" *) wire n3789_o;
  (* KEEP="TRUE" *) wire n3790_o;
  (* KEEP="TRUE" *) wire n3791_o;
  (* KEEP="TRUE" *) wire n3792_o;
  (* KEEP="TRUE" *) wire n3793_o;
  (* KEEP="TRUE" *) wire n3794_o;
  (* KEEP="TRUE" *) wire n3795_o;
  (* KEEP="TRUE" *) wire n3796_o;
  (* KEEP="TRUE" *) wire n3797_o;
  (* KEEP="TRUE" *) wire n3798_o;
  (* KEEP="TRUE" *) wire n3799_o;
  (* KEEP="TRUE" *) wire n3800_o;
  (* KEEP="TRUE" *) wire n3801_o;
  (* KEEP="TRUE" *) wire n3802_o;
  (* KEEP="TRUE" *) wire n3803_o;
  (* KEEP="TRUE" *) wire n3804_o;
  (* KEEP="TRUE" *) wire n3805_o;
  (* KEEP="TRUE" *) wire n3806_o;
  (* KEEP="TRUE" *) wire n3807_o;
  (* KEEP="TRUE" *) wire n3808_o;
  (* KEEP="TRUE" *) wire n3809_o;
  (* KEEP="TRUE" *) wire n3810_o;
  (* KEEP="TRUE" *) wire n3811_o;
  (* KEEP="TRUE" *) wire n3812_o;
  (* KEEP="TRUE" *) wire n3813_o;
  (* KEEP="TRUE" *) wire n3814_o;
  (* KEEP="TRUE" *) wire n3815_o;
  (* KEEP="TRUE" *) wire n3816_o;
  (* KEEP="TRUE" *) wire n3817_o;
  (* KEEP="TRUE" *) wire n3818_o;
  (* KEEP="TRUE" *) wire n3819_o;
  (* KEEP="TRUE" *) wire n3820_o;
  (* KEEP="TRUE" *) wire n3821_o;
  (* KEEP="TRUE" *) wire n3822_o;
  (* KEEP="TRUE" *) wire n3823_o;
  (* KEEP="TRUE" *) wire n3824_o;
  (* KEEP="TRUE" *) wire n3825_o;
  (* KEEP="TRUE" *) wire n3826_o;
  (* KEEP="TRUE" *) wire n3827_o;
  (* KEEP="TRUE" *) wire n3828_o;
  (* KEEP="TRUE" *) wire n3829_o;
  (* KEEP="TRUE" *) wire n3830_o;
  (* KEEP="TRUE" *) wire n3831_o;
  (* KEEP="TRUE" *) wire n3832_o;
  (* KEEP="TRUE" *) wire n3833_o;
  (* KEEP="TRUE" *) wire n3834_o;
  (* KEEP="TRUE" *) wire n3835_o;
  (* KEEP="TRUE" *) wire n3836_o;
  (* KEEP="TRUE" *) wire n3837_o;
  (* KEEP="TRUE" *) wire n3838_o;
  (* KEEP="TRUE" *) wire n3839_o;
  (* KEEP="TRUE" *) wire n3840_o;
  (* KEEP="TRUE" *) wire n3841_o;
  (* KEEP="TRUE" *) wire n3842_o;
  (* KEEP="TRUE" *) wire n3843_o;
  (* KEEP="TRUE" *) wire n3844_o;
  (* KEEP="TRUE" *) wire n3845_o;
  (* KEEP="TRUE" *) wire n3846_o;
  (* KEEP="TRUE" *) wire n3847_o;
  (* KEEP="TRUE" *) wire n3848_o;
  (* KEEP="TRUE" *) wire n3849_o;
  (* KEEP="TRUE" *) wire n3850_o;
  (* KEEP="TRUE" *) wire n3851_o;
  (* KEEP="TRUE" *) wire n3852_o;
  (* KEEP="TRUE" *) wire n3853_o;
  (* KEEP="TRUE" *) wire n3854_o;
  (* KEEP="TRUE" *) wire n3855_o;
  (* KEEP="TRUE" *) wire n3856_o;
  (* KEEP="TRUE" *) wire n3857_o;
  (* KEEP="TRUE" *) wire n3858_o;
  (* KEEP="TRUE" *) wire n3859_o;
  (* KEEP="TRUE" *) wire n3860_o;
  (* KEEP="TRUE" *) wire n3861_o;
  (* KEEP="TRUE" *) wire n3862_o;
  (* KEEP="TRUE" *) wire n3863_o;
  (* KEEP="TRUE" *) wire n3864_o;
  (* KEEP="TRUE" *) wire n3865_o;
  (* KEEP="TRUE" *) wire n3866_o;
  (* KEEP="TRUE" *) wire n3867_o;
  (* KEEP="TRUE" *) wire n3868_o;
  (* KEEP="TRUE" *) wire n3869_o;
  (* KEEP="TRUE" *) wire n3870_o;
  (* KEEP="TRUE" *) wire n3871_o;
  (* KEEP="TRUE" *) wire n3872_o;
  (* KEEP="TRUE" *) wire n3873_o;
  (* KEEP="TRUE" *) wire n3874_o;
  (* KEEP="TRUE" *) wire n3875_o;
  (* KEEP="TRUE" *) wire n3876_o;
  (* KEEP="TRUE" *) wire n3877_o;
  (* KEEP="TRUE" *) wire n3878_o;
  (* KEEP="TRUE" *) wire n3879_o;
  (* KEEP="TRUE" *) wire n3880_o;
  (* KEEP="TRUE" *) wire n3881_o;
  (* KEEP="TRUE" *) wire n3882_o;
  (* KEEP="TRUE" *) wire n3883_o;
  (* KEEP="TRUE" *) wire n3884_o;
  (* KEEP="TRUE" *) wire n3885_o;
  (* KEEP="TRUE" *) wire n3886_o;
  (* KEEP="TRUE" *) wire n3887_o;
  (* KEEP="TRUE" *) wire n3888_o;
  (* KEEP="TRUE" *) wire n3889_o;
  (* KEEP="TRUE" *) wire n3890_o;
  (* KEEP="TRUE" *) wire n3891_o;
  (* KEEP="TRUE" *) wire n3892_o;
  (* KEEP="TRUE" *) wire n3893_o;
  (* KEEP="TRUE" *) wire n3894_o;
  (* KEEP="TRUE" *) wire n3895_o;
  (* KEEP="TRUE" *) wire n3896_o;
  (* KEEP="TRUE" *) wire n3897_o;
  (* KEEP="TRUE" *) wire n3898_o;
  (* KEEP="TRUE" *) wire n3899_o;
  (* KEEP="TRUE" *) wire n3900_o;
  (* KEEP="TRUE" *) wire n3901_o;
  (* KEEP="TRUE" *) wire n3902_o;
  (* KEEP="TRUE" *) wire n3903_o;
  (* KEEP="TRUE" *) wire n3904_o;
  (* KEEP="TRUE" *) wire n3905_o;
  (* KEEP="TRUE" *) wire n3906_o;
  (* KEEP="TRUE" *) wire n3907_o;
  (* KEEP="TRUE" *) wire n3908_o;
  (* KEEP="TRUE" *) wire n3909_o;
  (* KEEP="TRUE" *) wire n3910_o;
  (* KEEP="TRUE" *) wire n3911_o;
  (* KEEP="TRUE" *) wire n3912_o;
  (* KEEP="TRUE" *) wire n3913_o;
  (* KEEP="TRUE" *) wire n3914_o;
  (* KEEP="TRUE" *) wire n3915_o;
  (* KEEP="TRUE" *) wire n3916_o;
  (* KEEP="TRUE" *) wire n3917_o;
  (* KEEP="TRUE" *) wire n3918_o;
  (* KEEP="TRUE" *) wire n3919_o;
  (* KEEP="TRUE" *) wire n3920_o;
  (* KEEP="TRUE" *) wire n3921_o;
  (* KEEP="TRUE" *) wire n3922_o;
  (* KEEP="TRUE" *) wire n3923_o;
  (* KEEP="TRUE" *) wire n3924_o;
  (* KEEP="TRUE" *) wire n3925_o;
  (* KEEP="TRUE" *) wire n3926_o;
  (* KEEP="TRUE" *) wire n3927_o;
  (* KEEP="TRUE" *) wire n3928_o;
  (* KEEP="TRUE" *) wire n3929_o;
  (* KEEP="TRUE" *) wire n3930_o;
  (* KEEP="TRUE" *) wire n3931_o;
  (* KEEP="TRUE" *) wire n3932_o;
  (* KEEP="TRUE" *) wire n3933_o;
  (* KEEP="TRUE" *) wire n3934_o;
  (* KEEP="TRUE" *) wire n3935_o;
  (* KEEP="TRUE" *) wire n3936_o;
  (* KEEP="TRUE" *) wire n3937_o;
  (* KEEP="TRUE" *) wire n3938_o;
  (* KEEP="TRUE" *) wire n3939_o;
  (* KEEP="TRUE" *) wire n3940_o;
  (* KEEP="TRUE" *) wire n3941_o;
  (* KEEP="TRUE" *) wire n3942_o;
  (* KEEP="TRUE" *) wire n3943_o;
  (* KEEP="TRUE" *) wire n3944_o;
  (* KEEP="TRUE" *) wire n3945_o;
  (* KEEP="TRUE" *) wire n3946_o;
  (* KEEP="TRUE" *) wire n3947_o;
  (* KEEP="TRUE" *) wire n3948_o;
  (* KEEP="TRUE" *) wire n3949_o;
  (* KEEP="TRUE" *) wire n3950_o;
  (* KEEP="TRUE" *) wire n3951_o;
  (* KEEP="TRUE" *) wire n3952_o;
  (* KEEP="TRUE" *) wire n3953_o;
  (* KEEP="TRUE" *) wire n3954_o;
  (* KEEP="TRUE" *) wire n3955_o;
  (* KEEP="TRUE" *) wire n3956_o;
  (* KEEP="TRUE" *) wire n3957_o;
  (* KEEP="TRUE" *) wire n3958_o;
  (* KEEP="TRUE" *) wire n3959_o;
  (* KEEP="TRUE" *) wire n3960_o;
  (* KEEP="TRUE" *) wire n3961_o;
  (* KEEP="TRUE" *) wire n3962_o;
  (* KEEP="TRUE" *) wire n3963_o;
  (* KEEP="TRUE" *) wire n3964_o;
  (* KEEP="TRUE" *) wire n3965_o;
  (* KEEP="TRUE" *) wire n3966_o;
  (* KEEP="TRUE" *) wire n3967_o;
  (* KEEP="TRUE" *) wire n3968_o;
  (* KEEP="TRUE" *) wire n3969_o;
  (* KEEP="TRUE" *) wire n3970_o;
  (* KEEP="TRUE" *) wire n3971_o;
  (* KEEP="TRUE" *) wire n3972_o;
  (* KEEP="TRUE" *) wire n3973_o;
  (* KEEP="TRUE" *) wire n3974_o;
  (* KEEP="TRUE" *) wire n3975_o;
  (* KEEP="TRUE" *) wire n3976_o;
  (* KEEP="TRUE" *) wire n3977_o;
  (* KEEP="TRUE" *) wire n3978_o;
  (* KEEP="TRUE" *) wire n3979_o;
  (* KEEP="TRUE" *) wire n3980_o;
  (* KEEP="TRUE" *) wire n3981_o;
  (* KEEP="TRUE" *) wire n3982_o;
  (* KEEP="TRUE" *) wire n3983_o;
  (* KEEP="TRUE" *) wire n3984_o;
  (* KEEP="TRUE" *) wire n3985_o;
  (* KEEP="TRUE" *) wire n3986_o;
  (* KEEP="TRUE" *) wire n3987_o;
  (* KEEP="TRUE" *) wire n3988_o;
  (* KEEP="TRUE" *) wire n3989_o;
  (* KEEP="TRUE" *) wire n3990_o;
  (* KEEP="TRUE" *) wire n3991_o;
  (* KEEP="TRUE" *) wire n3992_o;
  (* KEEP="TRUE" *) wire n3993_o;
  (* KEEP="TRUE" *) wire n3994_o;
  (* KEEP="TRUE" *) wire n3995_o;
  (* KEEP="TRUE" *) wire n3996_o;
  (* KEEP="TRUE" *) wire n3997_o;
  (* KEEP="TRUE" *) wire n3998_o;
  (* KEEP="TRUE" *) wire n3999_o;
  (* KEEP="TRUE" *) wire n4000_o;
  (* KEEP="TRUE" *) wire n4001_o;
  (* KEEP="TRUE" *) wire n4002_o;
  (* KEEP="TRUE" *) wire n4003_o;
  (* KEEP="TRUE" *) wire n4004_o;
  (* KEEP="TRUE" *) wire n4005_o;
  (* KEEP="TRUE" *) wire n4006_o;
  (* KEEP="TRUE" *) wire n4007_o;
  (* KEEP="TRUE" *) wire n4008_o;
  (* KEEP="TRUE" *) wire n4009_o;
  (* KEEP="TRUE" *) wire n4010_o;
  (* KEEP="TRUE" *) wire n4011_o;
  (* KEEP="TRUE" *) wire n4012_o;
  (* KEEP="TRUE" *) wire n4013_o;
  (* KEEP="TRUE" *) wire n4014_o;
  (* KEEP="TRUE" *) wire n4015_o;
  (* KEEP="TRUE" *) wire n4016_o;
  (* KEEP="TRUE" *) wire n4017_o;
  (* KEEP="TRUE" *) wire n4018_o;
  (* KEEP="TRUE" *) wire n4019_o;
  (* KEEP="TRUE" *) wire n4020_o;
  (* KEEP="TRUE" *) wire n4021_o;
  (* KEEP="TRUE" *) wire n4022_o;
  (* KEEP="TRUE" *) wire n4023_o;
  (* KEEP="TRUE" *) wire n4024_o;
  (* KEEP="TRUE" *) wire n4025_o;
  (* KEEP="TRUE" *) wire n4026_o;
  (* KEEP="TRUE" *) wire n4027_o;
  (* KEEP="TRUE" *) wire n4028_o;
  (* KEEP="TRUE" *) wire n4029_o;
  (* KEEP="TRUE" *) wire n4030_o;
  (* KEEP="TRUE" *) wire n4031_o;
  (* KEEP="TRUE" *) wire n4032_o;
  (* KEEP="TRUE" *) wire n4033_o;
  (* KEEP="TRUE" *) wire n4034_o;
  (* KEEP="TRUE" *) wire n4035_o;
  (* KEEP="TRUE" *) wire n4036_o;
  (* KEEP="TRUE" *) wire n4037_o;
  (* KEEP="TRUE" *) wire n4038_o;
  (* KEEP="TRUE" *) wire n4039_o;
  (* KEEP="TRUE" *) wire n4040_o;
  (* KEEP="TRUE" *) wire n4041_o;
  (* KEEP="TRUE" *) wire n4042_o;
  (* KEEP="TRUE" *) wire n4043_o;
  (* KEEP="TRUE" *) wire n4044_o;
  (* KEEP="TRUE" *) wire n4045_o;
  (* KEEP="TRUE" *) wire n4046_o;
  (* KEEP="TRUE" *) wire n4047_o;
  (* KEEP="TRUE" *) wire n4048_o;
  (* KEEP="TRUE" *) wire n4049_o;
  (* KEEP="TRUE" *) wire n4050_o;
  (* KEEP="TRUE" *) wire n4051_o;
  (* KEEP="TRUE" *) wire n4052_o;
  (* KEEP="TRUE" *) wire n4053_o;
  (* KEEP="TRUE" *) wire n4054_o;
  (* KEEP="TRUE" *) wire n4055_o;
  (* KEEP="TRUE" *) wire n4056_o;
  (* KEEP="TRUE" *) wire n4057_o;
  (* KEEP="TRUE" *) wire n4058_o;
  (* KEEP="TRUE" *) wire n4059_o;
  (* KEEP="TRUE" *) wire n4060_o;
  (* KEEP="TRUE" *) wire n4061_o;
  (* KEEP="TRUE" *) wire n4062_o;
  (* KEEP="TRUE" *) wire n4063_o;
  (* KEEP="TRUE" *) wire n4064_o;
  (* KEEP="TRUE" *) wire n4065_o;
  (* KEEP="TRUE" *) wire n4066_o;
  (* KEEP="TRUE" *) wire n4067_o;
  (* KEEP="TRUE" *) wire n4068_o;
  (* KEEP="TRUE" *) wire n4069_o;
  (* KEEP="TRUE" *) wire n4070_o;
  (* KEEP="TRUE" *) wire n4071_o;
  (* KEEP="TRUE" *) wire n4072_o;
  (* KEEP="TRUE" *) wire n4073_o;
  (* KEEP="TRUE" *) wire n4074_o;
  (* KEEP="TRUE" *) wire n4075_o;
  (* KEEP="TRUE" *) wire n4076_o;
  (* KEEP="TRUE" *) wire n4077_o;
  (* KEEP="TRUE" *) wire n4078_o;
  (* KEEP="TRUE" *) wire n4079_o;
  (* KEEP="TRUE" *) wire n4080_o;
  (* KEEP="TRUE" *) wire n4081_o;
  (* KEEP="TRUE" *) wire n4082_o;
  (* KEEP="TRUE" *) wire n4083_o;
  (* KEEP="TRUE" *) wire n4084_o;
  (* KEEP="TRUE" *) wire n4085_o;
  (* KEEP="TRUE" *) wire n4086_o;
  (* KEEP="TRUE" *) wire n4087_o;
  (* KEEP="TRUE" *) wire n4088_o;
  (* KEEP="TRUE" *) wire n4089_o;
  (* KEEP="TRUE" *) wire n4090_o;
  (* KEEP="TRUE" *) wire n4091_o;
  (* KEEP="TRUE" *) wire n4092_o;
  (* KEEP="TRUE" *) wire n4093_o;
  (* KEEP="TRUE" *) wire n4094_o;
  (* KEEP="TRUE" *) wire n4095_o;
  (* KEEP="TRUE" *) wire n4096_o;
  (* KEEP="TRUE" *) wire n4097_o;
  (* KEEP="TRUE" *) wire n4098_o;
  (* KEEP="TRUE" *) wire n4099_o;
  (* KEEP="TRUE" *) wire n4100_o;
  (* KEEP="TRUE" *) wire n4101_o;
  (* KEEP="TRUE" *) wire n4102_o;
  (* KEEP="TRUE" *) wire n4103_o;
  (* KEEP="TRUE" *) wire n4104_o;
  (* KEEP="TRUE" *) wire n4105_o;
  (* KEEP="TRUE" *) wire n4106_o;
  (* KEEP="TRUE" *) wire n4107_o;
  (* KEEP="TRUE" *) wire n4108_o;
  (* KEEP="TRUE" *) wire n4109_o;
  (* KEEP="TRUE" *) wire n4110_o;
  (* KEEP="TRUE" *) wire n4111_o;
  (* KEEP="TRUE" *) wire n4112_o;
  (* KEEP="TRUE" *) wire n4113_o;
  (* KEEP="TRUE" *) wire n4114_o;
  (* KEEP="TRUE" *) wire n4115_o;
  (* KEEP="TRUE" *) wire n4116_o;
  (* KEEP="TRUE" *) wire n4117_o;
  (* KEEP="TRUE" *) wire n4118_o;
  (* KEEP="TRUE" *) wire n4119_o;
  (* KEEP="TRUE" *) wire n4120_o;
  (* KEEP="TRUE" *) wire n4121_o;
  (* KEEP="TRUE" *) wire n4122_o;
  (* KEEP="TRUE" *) wire n4123_o;
  (* KEEP="TRUE" *) wire n4124_o;
  (* KEEP="TRUE" *) wire n4125_o;
  (* KEEP="TRUE" *) wire n4126_o;
  (* KEEP="TRUE" *) wire n4127_o;
  (* KEEP="TRUE" *) wire n4128_o;
  (* KEEP="TRUE" *) wire n4129_o;
  (* KEEP="TRUE" *) wire n4130_o;
  (* KEEP="TRUE" *) wire n4131_o;
  (* KEEP="TRUE" *) wire n4132_o;
  (* KEEP="TRUE" *) wire n4133_o;
  (* KEEP="TRUE" *) wire n4134_o;
  (* KEEP="TRUE" *) wire n4135_o;
  (* KEEP="TRUE" *) wire n4136_o;
  (* KEEP="TRUE" *) wire n4137_o;
  (* KEEP="TRUE" *) wire n4138_o;
  (* KEEP="TRUE" *) wire n4139_o;
  (* KEEP="TRUE" *) wire n4140_o;
  (* KEEP="TRUE" *) wire n4141_o;
  (* KEEP="TRUE" *) wire n4142_o;
  (* KEEP="TRUE" *) wire n4143_o;
  (* KEEP="TRUE" *) wire n4144_o;
  (* KEEP="TRUE" *) wire n4145_o;
  (* KEEP="TRUE" *) wire n4146_o;
  (* KEEP="TRUE" *) wire n4147_o;
  (* KEEP="TRUE" *) wire n4148_o;
  (* KEEP="TRUE" *) wire n4149_o;
  (* KEEP="TRUE" *) wire n4150_o;
  (* KEEP="TRUE" *) wire n4151_o;
  (* KEEP="TRUE" *) wire n4152_o;
  (* KEEP="TRUE" *) wire n4153_o;
  (* KEEP="TRUE" *) wire n4154_o;
  (* KEEP="TRUE" *) wire n4155_o;
  (* KEEP="TRUE" *) wire n4156_o;
  (* KEEP="TRUE" *) wire n4157_o;
  (* KEEP="TRUE" *) wire n4158_o;
  (* KEEP="TRUE" *) wire n4159_o;
  (* KEEP="TRUE" *) wire n4160_o;
  (* KEEP="TRUE" *) wire n4161_o;
  (* KEEP="TRUE" *) wire n4162_o;
  (* KEEP="TRUE" *) wire n4163_o;
  (* KEEP="TRUE" *) wire n4164_o;
  (* KEEP="TRUE" *) wire n4165_o;
  (* KEEP="TRUE" *) wire n4166_o;
  (* KEEP="TRUE" *) wire n4167_o;
  (* KEEP="TRUE" *) wire n4168_o;
  (* KEEP="TRUE" *) wire n4169_o;
  (* KEEP="TRUE" *) wire n4170_o;
  (* KEEP="TRUE" *) wire n4171_o;
  (* KEEP="TRUE" *) wire n4172_o;
  (* KEEP="TRUE" *) wire n4173_o;
  (* KEEP="TRUE" *) wire n4174_o;
  (* KEEP="TRUE" *) wire n4175_o;
  (* KEEP="TRUE" *) wire n4176_o;
  (* KEEP="TRUE" *) wire n4177_o;
  (* KEEP="TRUE" *) wire n4178_o;
  (* KEEP="TRUE" *) wire n4179_o;
  (* KEEP="TRUE" *) wire n4180_o;
  (* KEEP="TRUE" *) wire n4181_o;
  (* KEEP="TRUE" *) wire n4182_o;
  (* KEEP="TRUE" *) wire n4183_o;
  (* KEEP="TRUE" *) wire n4184_o;
  (* KEEP="TRUE" *) wire n4185_o;
  (* KEEP="TRUE" *) wire n4186_o;
  (* KEEP="TRUE" *) wire n4187_o;
  (* KEEP="TRUE" *) wire n4188_o;
  (* KEEP="TRUE" *) wire n4189_o;
  (* KEEP="TRUE" *) wire n4190_o;
  (* KEEP="TRUE" *) wire n4191_o;
  (* KEEP="TRUE" *) wire n4192_o;
  (* KEEP="TRUE" *) wire n4193_o;
  (* KEEP="TRUE" *) wire n4194_o;
  (* KEEP="TRUE" *) wire n4195_o;
  (* KEEP="TRUE" *) wire n4196_o;
  (* KEEP="TRUE" *) wire n4197_o;
  (* KEEP="TRUE" *) wire n4198_o;
  (* KEEP="TRUE" *) wire n4199_o;
  (* KEEP="TRUE" *) wire n4200_o;
  (* KEEP="TRUE" *) wire n4201_o;
  (* KEEP="TRUE" *) wire n4202_o;
  (* KEEP="TRUE" *) wire n4203_o;
  (* KEEP="TRUE" *) wire n4204_o;
  (* KEEP="TRUE" *) wire n4205_o;
  (* KEEP="TRUE" *) wire n4206_o;
  (* KEEP="TRUE" *) wire n4207_o;
  (* KEEP="TRUE" *) wire n4208_o;
  (* KEEP="TRUE" *) wire n4209_o;
  (* KEEP="TRUE" *) wire n4210_o;
  (* KEEP="TRUE" *) wire n4211_o;
  (* KEEP="TRUE" *) wire n4212_o;
  (* KEEP="TRUE" *) wire n4213_o;
  (* KEEP="TRUE" *) wire n4214_o;
  (* KEEP="TRUE" *) wire n4215_o;
  (* KEEP="TRUE" *) wire n4216_o;
  (* KEEP="TRUE" *) wire n4217_o;
  (* KEEP="TRUE" *) wire n4218_o;
  (* KEEP="TRUE" *) wire n4219_o;
  (* KEEP="TRUE" *) wire n4220_o;
  (* KEEP="TRUE" *) wire n4221_o;
  (* KEEP="TRUE" *) wire n4222_o;
  (* KEEP="TRUE" *) wire n4223_o;
  (* KEEP="TRUE" *) wire n4224_o;
  (* KEEP="TRUE" *) wire n4225_o;
  (* KEEP="TRUE" *) wire n4226_o;
  (* KEEP="TRUE" *) wire n4227_o;
  (* KEEP="TRUE" *) wire n4228_o;
  (* KEEP="TRUE" *) wire n4229_o;
  (* KEEP="TRUE" *) wire n4230_o;
  (* KEEP="TRUE" *) wire n4231_o;
  (* KEEP="TRUE" *) wire n4232_o;
  (* KEEP="TRUE" *) wire n4233_o;
  (* KEEP="TRUE" *) wire n4234_o;
  (* KEEP="TRUE" *) wire n4235_o;
  (* KEEP="TRUE" *) wire n4236_o;
  (* KEEP="TRUE" *) wire n4237_o;
  (* KEEP="TRUE" *) wire n4238_o;
  (* KEEP="TRUE" *) wire n4239_o;
  (* KEEP="TRUE" *) wire n4240_o;
  (* KEEP="TRUE" *) wire n4241_o;
  (* KEEP="TRUE" *) wire n4242_o;
  (* KEEP="TRUE" *) wire n4243_o;
  (* KEEP="TRUE" *) wire n4244_o;
  (* KEEP="TRUE" *) wire n4245_o;
  (* KEEP="TRUE" *) wire n4246_o;
  (* KEEP="TRUE" *) wire n4247_o;
  (* KEEP="TRUE" *) wire n4248_o;
  (* KEEP="TRUE" *) wire n4249_o;
  (* KEEP="TRUE" *) wire n4250_o;
  (* KEEP="TRUE" *) wire n4251_o;
  (* KEEP="TRUE" *) wire n4252_o;
  (* KEEP="TRUE" *) wire n4253_o;
  (* KEEP="TRUE" *) wire n4254_o;
  (* KEEP="TRUE" *) wire n4255_o;
  (* KEEP="TRUE" *) wire n4256_o;
  (* KEEP="TRUE" *) wire n4257_o;
  (* KEEP="TRUE" *) wire n4258_o;
  (* KEEP="TRUE" *) wire n4259_o;
  (* KEEP="TRUE" *) wire n4260_o;
  (* KEEP="TRUE" *) wire n4261_o;
  (* KEEP="TRUE" *) wire n4262_o;
  (* KEEP="TRUE" *) wire n4263_o;
  (* KEEP="TRUE" *) wire n4264_o;
  (* KEEP="TRUE" *) wire n4265_o;
  (* KEEP="TRUE" *) wire n4266_o;
  (* KEEP="TRUE" *) wire n4267_o;
  (* KEEP="TRUE" *) wire n4268_o;
  (* KEEP="TRUE" *) wire n4269_o;
  (* KEEP="TRUE" *) wire n4270_o;
  (* KEEP="TRUE" *) wire n4271_o;
  (* KEEP="TRUE" *) wire n4272_o;
  (* KEEP="TRUE" *) wire n4273_o;
  (* KEEP="TRUE" *) wire n4274_o;
  (* KEEP="TRUE" *) wire n4275_o;
  (* KEEP="TRUE" *) wire n4276_o;
  (* KEEP="TRUE" *) wire n4277_o;
  (* KEEP="TRUE" *) wire n4278_o;
  (* KEEP="TRUE" *) wire n4279_o;
  (* KEEP="TRUE" *) wire n4280_o;
  (* KEEP="TRUE" *) wire n4281_o;
  (* KEEP="TRUE" *) wire n4282_o;
  (* KEEP="TRUE" *) wire n4283_o;
  (* KEEP="TRUE" *) wire n4284_o;
  (* KEEP="TRUE" *) wire n4285_o;
  (* KEEP="TRUE" *) wire n4286_o;
  (* KEEP="TRUE" *) wire n4287_o;
  (* KEEP="TRUE" *) wire n4288_o;
  (* KEEP="TRUE" *) wire n4289_o;
  (* KEEP="TRUE" *) wire n4290_o;
  (* KEEP="TRUE" *) wire n4291_o;
  (* KEEP="TRUE" *) wire n4292_o;
  (* KEEP="TRUE" *) wire n4293_o;
  (* KEEP="TRUE" *) wire n4294_o;
  (* KEEP="TRUE" *) wire n4295_o;
  (* KEEP="TRUE" *) wire n4296_o;
  (* KEEP="TRUE" *) wire n4297_o;
  (* KEEP="TRUE" *) wire n4298_o;
  (* KEEP="TRUE" *) wire n4299_o;
  (* KEEP="TRUE" *) wire n4300_o;
  (* KEEP="TRUE" *) wire n4301_o;
  (* KEEP="TRUE" *) wire n4302_o;
  (* KEEP="TRUE" *) wire n4303_o;
  (* KEEP="TRUE" *) wire n4304_o;
  (* KEEP="TRUE" *) wire n4305_o;
  (* KEEP="TRUE" *) wire n4306_o;
  (* KEEP="TRUE" *) wire n4307_o;
  (* KEEP="TRUE" *) wire n4308_o;
  (* KEEP="TRUE" *) wire n4309_o;
  (* KEEP="TRUE" *) wire n4310_o;
  (* KEEP="TRUE" *) wire n4311_o;
  (* KEEP="TRUE" *) wire n4312_o;
  (* KEEP="TRUE" *) wire n4313_o;
  (* KEEP="TRUE" *) wire n4314_o;
  (* KEEP="TRUE" *) wire n4315_o;
  (* KEEP="TRUE" *) wire n4316_o;
  (* KEEP="TRUE" *) wire n4317_o;
  (* KEEP="TRUE" *) wire n4318_o;
  (* KEEP="TRUE" *) wire n4319_o;
  (* KEEP="TRUE" *) wire n4320_o;
  (* KEEP="TRUE" *) wire n4321_o;
  (* KEEP="TRUE" *) wire n4322_o;
  (* KEEP="TRUE" *) wire n4323_o;
  (* KEEP="TRUE" *) wire n4324_o;
  (* KEEP="TRUE" *) wire n4325_o;
  (* KEEP="TRUE" *) wire n4326_o;
  (* KEEP="TRUE" *) wire n4327_o;
  (* KEEP="TRUE" *) wire n4328_o;
  (* KEEP="TRUE" *) wire n4329_o;
  (* KEEP="TRUE" *) wire n4330_o;
  (* KEEP="TRUE" *) wire n4331_o;
  (* KEEP="TRUE" *) wire n4332_o;
  (* KEEP="TRUE" *) wire n4333_o;
  (* KEEP="TRUE" *) wire n4334_o;
  (* KEEP="TRUE" *) wire n4335_o;
  (* KEEP="TRUE" *) wire n4336_o;
  (* KEEP="TRUE" *) wire n4337_o;
  (* KEEP="TRUE" *) wire n4338_o;
  (* KEEP="TRUE" *) wire n4339_o;
  (* KEEP="TRUE" *) wire n4340_o;
  (* KEEP="TRUE" *) wire n4341_o;
  (* KEEP="TRUE" *) wire n4342_o;
  (* KEEP="TRUE" *) wire n4343_o;
  (* KEEP="TRUE" *) wire n4344_o;
  (* KEEP="TRUE" *) wire n4345_o;
  (* KEEP="TRUE" *) wire n4346_o;
  (* KEEP="TRUE" *) wire n4347_o;
  (* KEEP="TRUE" *) wire n4348_o;
  (* KEEP="TRUE" *) wire n4349_o;
  (* KEEP="TRUE" *) wire n4350_o;
  (* KEEP="TRUE" *) wire n4351_o;
  (* KEEP="TRUE" *) wire n4352_o;
  (* KEEP="TRUE" *) wire n4353_o;
  (* KEEP="TRUE" *) wire n4354_o;
  (* KEEP="TRUE" *) wire n4355_o;
  (* KEEP="TRUE" *) wire n4356_o;
  (* KEEP="TRUE" *) wire n4357_o;
  (* KEEP="TRUE" *) wire n4358_o;
  (* KEEP="TRUE" *) wire n4359_o;
  (* KEEP="TRUE" *) wire n4360_o;
  (* KEEP="TRUE" *) wire n4361_o;
  (* KEEP="TRUE" *) wire n4362_o;
  (* KEEP="TRUE" *) wire n4363_o;
  (* KEEP="TRUE" *) wire n4364_o;
  (* KEEP="TRUE" *) wire n4365_o;
  (* KEEP="TRUE" *) wire n4366_o;
  (* KEEP="TRUE" *) wire n4367_o;
  (* KEEP="TRUE" *) wire n4368_o;
  (* KEEP="TRUE" *) wire n4369_o;
  (* KEEP="TRUE" *) wire n4370_o;
  (* KEEP="TRUE" *) wire n4371_o;
  (* KEEP="TRUE" *) wire n4372_o;
  (* KEEP="TRUE" *) wire n4373_o;
  (* KEEP="TRUE" *) wire n4374_o;
  (* KEEP="TRUE" *) wire n4375_o;
  (* KEEP="TRUE" *) wire n4376_o;
  (* KEEP="TRUE" *) wire n4377_o;
  (* KEEP="TRUE" *) wire n4378_o;
  (* KEEP="TRUE" *) wire n4379_o;
  (* KEEP="TRUE" *) wire n4380_o;
  (* KEEP="TRUE" *) wire n4381_o;
  (* KEEP="TRUE" *) wire n4382_o;
  (* KEEP="TRUE" *) wire n4383_o;
  (* KEEP="TRUE" *) wire n4384_o;
  (* KEEP="TRUE" *) wire n4385_o;
  (* KEEP="TRUE" *) wire n4386_o;
  (* KEEP="TRUE" *) wire n4387_o;
  (* KEEP="TRUE" *) wire n4388_o;
  (* KEEP="TRUE" *) wire n4389_o;
  (* KEEP="TRUE" *) wire n4390_o;
  (* KEEP="TRUE" *) wire n4391_o;
  (* KEEP="TRUE" *) wire n4392_o;
  (* KEEP="TRUE" *) wire n4393_o;
  (* KEEP="TRUE" *) wire n4394_o;
  (* KEEP="TRUE" *) wire n4395_o;
  (* KEEP="TRUE" *) wire n4396_o;
  (* KEEP="TRUE" *) wire n4397_o;
  (* KEEP="TRUE" *) wire n4398_o;
  (* KEEP="TRUE" *) wire n4399_o;
  (* KEEP="TRUE" *) wire n4400_o;
  (* KEEP="TRUE" *) wire n4401_o;
  (* KEEP="TRUE" *) wire n4402_o;
  (* KEEP="TRUE" *) wire n4403_o;
  (* KEEP="TRUE" *) wire n4404_o;
  (* KEEP="TRUE" *) wire n4405_o;
  (* KEEP="TRUE" *) wire n4406_o;
  (* KEEP="TRUE" *) wire n4407_o;
  (* KEEP="TRUE" *) wire n4408_o;
  (* KEEP="TRUE" *) wire n4409_o;
  (* KEEP="TRUE" *) wire n4410_o;
  (* KEEP="TRUE" *) wire n4411_o;
  (* KEEP="TRUE" *) wire n4412_o;
  (* KEEP="TRUE" *) wire n4413_o;
  (* KEEP="TRUE" *) wire n4414_o;
  (* KEEP="TRUE" *) wire n4415_o;
  (* KEEP="TRUE" *) wire n4416_o;
  (* KEEP="TRUE" *) wire n4417_o;
  (* KEEP="TRUE" *) wire n4418_o;
  (* KEEP="TRUE" *) wire n4419_o;
  (* KEEP="TRUE" *) wire n4420_o;
  (* KEEP="TRUE" *) wire n4421_o;
  (* KEEP="TRUE" *) wire n4422_o;
  (* KEEP="TRUE" *) wire n4423_o;
  (* KEEP="TRUE" *) wire n4424_o;
  (* KEEP="TRUE" *) wire n4425_o;
  (* KEEP="TRUE" *) wire n4426_o;
  (* KEEP="TRUE" *) wire n4427_o;
  (* KEEP="TRUE" *) wire n4428_o;
  (* KEEP="TRUE" *) wire n4429_o;
  (* KEEP="TRUE" *) wire n4430_o;
  (* KEEP="TRUE" *) wire n4431_o;
  (* KEEP="TRUE" *) wire n4432_o;
  (* KEEP="TRUE" *) wire n4433_o;
  (* KEEP="TRUE" *) wire n4434_o;
  (* KEEP="TRUE" *) wire n4435_o;
  (* KEEP="TRUE" *) wire n4436_o;
  (* KEEP="TRUE" *) wire n4437_o;
  (* KEEP="TRUE" *) wire n4438_o;
  (* KEEP="TRUE" *) wire n4439_o;
  (* KEEP="TRUE" *) wire n4440_o;
  (* KEEP="TRUE" *) wire n4441_o;
  (* KEEP="TRUE" *) wire n4442_o;
  (* KEEP="TRUE" *) wire n4443_o;
  (* KEEP="TRUE" *) wire n4444_o;
  (* KEEP="TRUE" *) wire n4445_o;
  (* KEEP="TRUE" *) wire n4446_o;
  (* KEEP="TRUE" *) wire n4447_o;
  (* KEEP="TRUE" *) wire n4448_o;
  (* KEEP="TRUE" *) wire n4449_o;
  (* KEEP="TRUE" *) wire n4450_o;
  (* KEEP="TRUE" *) wire n4451_o;
  (* KEEP="TRUE" *) wire n4452_o;
  (* KEEP="TRUE" *) wire n4453_o;
  (* KEEP="TRUE" *) wire n4454_o;
  (* KEEP="TRUE" *) wire n4455_o;
  (* KEEP="TRUE" *) wire n4456_o;
  (* KEEP="TRUE" *) wire n4457_o;
  (* KEEP="TRUE" *) wire n4458_o;
  (* KEEP="TRUE" *) wire n4459_o;
  (* KEEP="TRUE" *) wire n4460_o;
  (* KEEP="TRUE" *) wire n4461_o;
  (* KEEP="TRUE" *) wire n4462_o;
  (* KEEP="TRUE" *) wire n4463_o;
  (* KEEP="TRUE" *) wire n4464_o;
  (* KEEP="TRUE" *) wire n4465_o;
  (* KEEP="TRUE" *) wire n4466_o;
  (* KEEP="TRUE" *) wire n4467_o;
  (* KEEP="TRUE" *) wire n4468_o;
  (* KEEP="TRUE" *) wire n4469_o;
  (* KEEP="TRUE" *) wire n4470_o;
  (* KEEP="TRUE" *) wire n4471_o;
  (* KEEP="TRUE" *) wire n4472_o;
  (* KEEP="TRUE" *) wire n4473_o;
  (* KEEP="TRUE" *) wire n4474_o;
  (* KEEP="TRUE" *) wire n4475_o;
  (* KEEP="TRUE" *) wire n4476_o;
  (* KEEP="TRUE" *) wire n4477_o;
  (* KEEP="TRUE" *) wire n4478_o;
  (* KEEP="TRUE" *) wire n4479_o;
  (* KEEP="TRUE" *) wire n4480_o;
  (* KEEP="TRUE" *) wire n4481_o;
  (* KEEP="TRUE" *) wire n4482_o;
  (* KEEP="TRUE" *) wire n4483_o;
  (* KEEP="TRUE" *) wire n4484_o;
  (* KEEP="TRUE" *) wire n4485_o;
  (* KEEP="TRUE" *) wire n4486_o;
  (* KEEP="TRUE" *) wire n4487_o;
  (* KEEP="TRUE" *) wire n4488_o;
  (* KEEP="TRUE" *) wire n4489_o;
  (* KEEP="TRUE" *) wire n4490_o;
  (* KEEP="TRUE" *) wire n4491_o;
  (* KEEP="TRUE" *) wire n4492_o;
  (* KEEP="TRUE" *) wire n4493_o;
  (* KEEP="TRUE" *) wire n4494_o;
  (* KEEP="TRUE" *) wire n4495_o;
  (* KEEP="TRUE" *) wire n4496_o;
  (* KEEP="TRUE" *) wire n4497_o;
  (* KEEP="TRUE" *) wire n4498_o;
  (* KEEP="TRUE" *) wire n4499_o;
  (* KEEP="TRUE" *) wire n4500_o;
  (* KEEP="TRUE" *) wire n4501_o;
  (* KEEP="TRUE" *) wire n4502_o;
  (* KEEP="TRUE" *) wire n4503_o;
  (* KEEP="TRUE" *) wire n4504_o;
  (* KEEP="TRUE" *) wire n4505_o;
  (* KEEP="TRUE" *) wire n4506_o;
  (* KEEP="TRUE" *) wire n4507_o;
  (* KEEP="TRUE" *) wire n4508_o;
  (* KEEP="TRUE" *) wire n4509_o;
  (* KEEP="TRUE" *) wire n4510_o;
  (* KEEP="TRUE" *) wire n4511_o;
  (* KEEP="TRUE" *) wire n4512_o;
  (* KEEP="TRUE" *) wire n4513_o;
  (* KEEP="TRUE" *) wire n4514_o;
  (* KEEP="TRUE" *) wire n4515_o;
  (* KEEP="TRUE" *) wire n4516_o;
  (* KEEP="TRUE" *) wire n4517_o;
  (* KEEP="TRUE" *) wire n4518_o;
  (* KEEP="TRUE" *) wire n4519_o;
  (* KEEP="TRUE" *) wire n4520_o;
  (* KEEP="TRUE" *) wire n4521_o;
  (* KEEP="TRUE" *) wire n4522_o;
  (* KEEP="TRUE" *) wire n4523_o;
  (* KEEP="TRUE" *) wire n4524_o;
  (* KEEP="TRUE" *) wire n4525_o;
  (* KEEP="TRUE" *) wire n4526_o;
  (* KEEP="TRUE" *) wire n4527_o;
  (* KEEP="TRUE" *) wire n4528_o;
  (* KEEP="TRUE" *) wire n4529_o;
  (* KEEP="TRUE" *) wire n4530_o;
  (* KEEP="TRUE" *) wire n4531_o;
  (* KEEP="TRUE" *) wire n4532_o;
  (* KEEP="TRUE" *) wire n4533_o;
  (* KEEP="TRUE" *) wire n4534_o;
  (* KEEP="TRUE" *) wire n4535_o;
  (* KEEP="TRUE" *) wire n4536_o;
  (* KEEP="TRUE" *) wire n4537_o;
  (* KEEP="TRUE" *) wire n4538_o;
  (* KEEP="TRUE" *) wire n4539_o;
  (* KEEP="TRUE" *) wire n4540_o;
  (* KEEP="TRUE" *) wire n4541_o;
  (* KEEP="TRUE" *) wire n4542_o;
  (* KEEP="TRUE" *) wire n4543_o;
  (* KEEP="TRUE" *) wire n4544_o;
  (* KEEP="TRUE" *) wire n4545_o;
  (* KEEP="TRUE" *) wire n4546_o;
  (* KEEP="TRUE" *) wire n4547_o;
  (* KEEP="TRUE" *) wire n4548_o;
  (* KEEP="TRUE" *) wire n4549_o;
  (* KEEP="TRUE" *) wire n4550_o;
  (* KEEP="TRUE" *) wire n4551_o;
  (* KEEP="TRUE" *) wire n4552_o;
  (* KEEP="TRUE" *) wire n4553_o;
  (* KEEP="TRUE" *) wire n4554_o;
  (* KEEP="TRUE" *) wire n4555_o;
  (* KEEP="TRUE" *) wire n4556_o;
  (* KEEP="TRUE" *) wire n4557_o;
  (* KEEP="TRUE" *) wire n4558_o;
  (* KEEP="TRUE" *) wire n4559_o;
  (* KEEP="TRUE" *) wire n4560_o;
  (* KEEP="TRUE" *) wire n4561_o;
  (* KEEP="TRUE" *) wire n4562_o;
  (* KEEP="TRUE" *) wire n4563_o;
  (* KEEP="TRUE" *) wire n4564_o;
  (* KEEP="TRUE" *) wire n4565_o;
  (* KEEP="TRUE" *) wire n4566_o;
  (* KEEP="TRUE" *) wire n4567_o;
  (* KEEP="TRUE" *) wire n4568_o;
  (* KEEP="TRUE" *) wire n4569_o;
  (* KEEP="TRUE" *) wire n4570_o;
  (* KEEP="TRUE" *) wire n4571_o;
  (* KEEP="TRUE" *) wire n4572_o;
  (* KEEP="TRUE" *) wire n4573_o;
  (* KEEP="TRUE" *) wire n4574_o;
  (* KEEP="TRUE" *) wire n4575_o;
  (* KEEP="TRUE" *) wire n4576_o;
  (* KEEP="TRUE" *) wire n4577_o;
  (* KEEP="TRUE" *) wire n4578_o;
  (* KEEP="TRUE" *) wire n4579_o;
  (* KEEP="TRUE" *) wire n4580_o;
  (* KEEP="TRUE" *) wire n4581_o;
  (* KEEP="TRUE" *) wire n4582_o;
  (* KEEP="TRUE" *) wire n4583_o;
  (* KEEP="TRUE" *) wire n4584_o;
  (* KEEP="TRUE" *) wire n4585_o;
  (* KEEP="TRUE" *) wire n4586_o;
  (* KEEP="TRUE" *) wire n4587_o;
  (* KEEP="TRUE" *) wire n4588_o;
  (* KEEP="TRUE" *) wire n4589_o;
  (* KEEP="TRUE" *) wire n4590_o;
  (* KEEP="TRUE" *) wire n4591_o;
  (* KEEP="TRUE" *) wire n4592_o;
  (* KEEP="TRUE" *) wire n4593_o;
  (* KEEP="TRUE" *) wire n4594_o;
  (* KEEP="TRUE" *) wire n4595_o;
  (* KEEP="TRUE" *) wire n4596_o;
  (* KEEP="TRUE" *) wire n4597_o;
  (* KEEP="TRUE" *) wire n4598_o;
  (* KEEP="TRUE" *) wire n4599_o;
  (* KEEP="TRUE" *) wire n4600_o;
  (* KEEP="TRUE" *) wire n4601_o;
  (* KEEP="TRUE" *) wire n4602_o;
  (* KEEP="TRUE" *) wire n4603_o;
  (* KEEP="TRUE" *) wire n4604_o;
  (* KEEP="TRUE" *) wire n4605_o;
  (* KEEP="TRUE" *) wire n4606_o;
  (* KEEP="TRUE" *) wire n4607_o;
  (* KEEP="TRUE" *) wire n4608_o;
  (* KEEP="TRUE" *) wire n4609_o;
  (* KEEP="TRUE" *) wire n4610_o;
  (* KEEP="TRUE" *) wire n4611_o;
  (* KEEP="TRUE" *) wire n4612_o;
  (* KEEP="TRUE" *) wire n4613_o;
  (* KEEP="TRUE" *) wire n4614_o;
  (* KEEP="TRUE" *) wire n4615_o;
  (* KEEP="TRUE" *) wire n4616_o;
  (* KEEP="TRUE" *) wire n4617_o;
  (* KEEP="TRUE" *) wire n4618_o;
  (* KEEP="TRUE" *) wire n4619_o;
  (* KEEP="TRUE" *) wire n4620_o;
  (* KEEP="TRUE" *) wire n4621_o;
  (* KEEP="TRUE" *) wire n4622_o;
  (* KEEP="TRUE" *) wire n4623_o;
  (* KEEP="TRUE" *) wire n4624_o;
  (* KEEP="TRUE" *) wire n4625_o;
  (* KEEP="TRUE" *) wire n4626_o;
  (* KEEP="TRUE" *) wire n4627_o;
  (* KEEP="TRUE" *) wire n4628_o;
  (* KEEP="TRUE" *) wire n4629_o;
  (* KEEP="TRUE" *) wire n4630_o;
  (* KEEP="TRUE" *) wire n4631_o;
  (* KEEP="TRUE" *) wire n4632_o;
  (* KEEP="TRUE" *) wire n4633_o;
  (* KEEP="TRUE" *) wire n4634_o;
  (* KEEP="TRUE" *) wire n4635_o;
  (* KEEP="TRUE" *) wire n4636_o;
  (* KEEP="TRUE" *) wire n4637_o;
  (* KEEP="TRUE" *) wire n4638_o;
  (* KEEP="TRUE" *) wire n4639_o;
  (* KEEP="TRUE" *) wire n4640_o;
  (* KEEP="TRUE" *) wire n4641_o;
  (* KEEP="TRUE" *) wire n4642_o;
  (* KEEP="TRUE" *) wire n4643_o;
  (* KEEP="TRUE" *) wire [255:0] n4644_o;
  assign led1 = n487_q;
  assign led2 = n488_q;
  assign led3 = n187_o;
  assign led4 = n188_o;
  assign uart_tx = uart_tx_inst_tx_out;
  assign ledR_1 = n489_q;
  assign ledG_1 = n490_q;
  assign ledB_1 = n491_q;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:45:8  */
  assign received_word = uart_rx_inst_data_out; // (signal)
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:46:8  */
  assign rdy = uart_rx_inst_rdy; // (signal)
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:49:8  */
  always @*
    tx_en = n452_q; // (isignal)
  initial
    tx_en = 1'b0;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:50:8  */
  assign tx_busy = uart_tx_inst_busy_out; // (signal)
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:51:8  */
  always @*
    tx_data_in = n454_q; // (isignal)
  initial
    tx_data_in = 8'b00000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:55:8  */
  always @*
    shift_state = n455_q; // (isignal)
  initial
    shift_state = 1'b0;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:56:8  */
  always @*
    output_data = n456_q; // (isignal)
  initial
    output_data = 8'b00000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:106:8  */
  always @*
    internal_challenge_mux = n457_q; // (isignal)
  initial
    internal_challenge_mux = 8'b00000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:107:8  */
  always @*
    puf_response = n467_o; // (isignal)
  initial
    puf_response = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:108:8  */
  always @*
    puf_start = n184_o; // (isignal)
  initial
    puf_start = 1'b0;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:109:8  */
  always @*
    mux_1_challenge = n468_q; // (isignal)
  initial
    mux_1_challenge = 8'b00000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:110:8  */
  always @*
    mux_2_challenge = n469_q; // (isignal)
  initial
    mux_2_challenge = 8'b00000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:111:8  */
  always @*
    mux_1_out = uut1_n189; // (isignal)
  initial
    mux_1_out = 1'b0;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:112:8  */
  always @*
    mux_2_out = uut2_n192; // (isignal)
  initial
    mux_2_out = 1'b0;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:113:8  */
  always @*
    compteur_cycles = n470_q; // (isignal)
  initial
    compteur_cycles = 29'b00000000000000000000000000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:114:8  */
  always @*
    mux_1_counter = n472_q; // (isignal)
  initial
    mux_1_counter = 31'b0000000000000000000000000000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:115:8  */
  always @*
    mux_2_counter = n474_q; // (isignal)
  initial
    mux_2_counter = 31'b0000000000000000000000000000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:117:8  */
  always @*
    enable_1 = n475_q; // (isignal)
  initial
    enable_1 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:118:8  */
  always @*
    enable_2 = n476_q; // (isignal)
  initial
    enable_2 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:119:8  */
  always @*
    reset_counter = n477_q; // (isignal)
  initial
    reset_counter = 1'b0;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:120:8  */
  always @*
    enable_comparison = n478_q; // (isignal)
  initial
    enable_comparison = 1'b0;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:121:8  */
  always @*
    enable_counter = n479_q; // (isignal)
  initial
    enable_counter = 1'b0;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:123:8  */
  always @*
    data_valid = n480_q; // (isignal)
  initial
    data_valid = 1'b1;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:124:8  */
  always @*
    tx_available = n482_q; // (isignal)
  initial
    tx_available = 1'b1;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:125:8  */
  assign counter_timer = n186_o; // (signal)
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:126:8  */
  always @*
    timer_size = n216_o; // (isignal)
  initial
    timer_size = 32'b00000000000000000000000000000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:128:8  */
  always @*
    ro_filter = 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111; // (isignal)
  initial
    ro_filter = 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:129:8  */
  always @*
    rom_address = n483_q; // (isignal)
  initial
    rom_address = 8'b00000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:130:8  */
  assign rom_data_out = rom_n195; // (signal)
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:131:8  */
  always @*
    mode_select = n185_o; // (isignal)
  initial
    mode_select = 1'b0;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:135:8  */
  assign state = n484_q; // (signal)
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:138:8  */
  always @*
    transmission_state = n486_q; // (isignal)
  initial
    transmission_state = 5'b00000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:150:1  */
  uart_rx uart_rx_inst (
    .clk(clk),
    .rx_in(uart_rx),
    .busy_out(),
    .rdy(uart_rx_inst_rdy),
    .data_out(uart_rx_inst_data_out));
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:159:1  */
  uart_tx uart_tx_inst (
    .clk(clk),
    .reset(reset_btn),
    .data_in(tx_data_in),
    .en(tx_en),
    .busy_out(uart_tx_inst_busy_out),
    .tx_out(uart_tx_inst_tx_out));
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:172:20  */
  assign n47_o = ~tx_busy;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:178:21  */
  assign n50_o = data_valid ? 5'b00001 : 5'b00000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:175:17  */
  assign n52_o = transmission_state == 5'b00000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:186:56  */
  assign n53_o = puf_response[63:56];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:183:17  */
  assign n55_o = transmission_state == 5'b00001;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:188:17  */
  assign n57_o = transmission_state == 5'b00010;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:193:56  */
  assign n58_o = puf_response[55:48];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:191:17  */
  assign n60_o = transmission_state == 5'b00011;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:195:17  */
  assign n62_o = transmission_state == 5'b00100;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:200:56  */
  assign n63_o = puf_response[47:40];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:198:17  */
  assign n65_o = transmission_state == 5'b00101;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:202:17  */
  assign n67_o = transmission_state == 5'b00110;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:207:56  */
  assign n68_o = puf_response[39:32];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:205:17  */
  assign n70_o = transmission_state == 5'b00111;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:209:17  */
  assign n72_o = transmission_state == 5'b01000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:214:56  */
  assign n73_o = puf_response[31:24];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:212:17  */
  assign n75_o = transmission_state == 5'b01001;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:216:17  */
  assign n77_o = transmission_state == 5'b01010;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:221:56  */
  assign n78_o = puf_response[23:16];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:219:17  */
  assign n80_o = transmission_state == 5'b01011;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:223:17  */
  assign n82_o = transmission_state == 5'b01100;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:228:56  */
  assign n83_o = puf_response[15:8];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:226:17  */
  assign n85_o = transmission_state == 5'b01101;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:230:17  */
  assign n87_o = transmission_state == 5'b01110;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:235:56  */
  assign n88_o = puf_response[7:0];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:233:17  */
  assign n90_o = transmission_state == 5'b01111;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:237:25  */
  assign n92_o = transmission_state == 5'b10000;
  assign n93_o = {n92_o, n90_o, n87_o, n85_o, n82_o, n80_o, n77_o, n75_o, n72_o, n70_o, n67_o, n65_o, n62_o, n60_o, n57_o, n55_o, n52_o};
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:173:13  */
  always @*
    case (n93_o)
      17'b10000000000000000: n111_o = 1'b0;
      17'b01000000000000000: n111_o = 1'b1;
      17'b00100000000000000: n111_o = 1'b0;
      17'b00010000000000000: n111_o = 1'b1;
      17'b00001000000000000: n111_o = 1'b0;
      17'b00000100000000000: n111_o = 1'b1;
      17'b00000010000000000: n111_o = 1'b0;
      17'b00000001000000000: n111_o = 1'b1;
      17'b00000000100000000: n111_o = 1'b0;
      17'b00000000010000000: n111_o = 1'b1;
      17'b00000000001000000: n111_o = 1'b0;
      17'b00000000000100000: n111_o = 1'b1;
      17'b00000000000010000: n111_o = 1'b0;
      17'b00000000000001000: n111_o = 1'b1;
      17'b00000000000000100: n111_o = 1'b0;
      17'b00000000000000010: n111_o = 1'b1;
      17'b00000000000000001: n111_o = 1'b0;
      default: n111_o = tx_en;
    endcase
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:173:13  */
  always @*
    case (n93_o)
      17'b10000000000000000: n112_o = tx_data_in;
      17'b01000000000000000: n112_o = n88_o;
      17'b00100000000000000: n112_o = tx_data_in;
      17'b00010000000000000: n112_o = n83_o;
      17'b00001000000000000: n112_o = tx_data_in;
      17'b00000100000000000: n112_o = n78_o;
      17'b00000010000000000: n112_o = tx_data_in;
      17'b00000001000000000: n112_o = n73_o;
      17'b00000000100000000: n112_o = tx_data_in;
      17'b00000000010000000: n112_o = n68_o;
      17'b00000000001000000: n112_o = tx_data_in;
      17'b00000000000100000: n112_o = n63_o;
      17'b00000000000010000: n112_o = tx_data_in;
      17'b00000000000001000: n112_o = n58_o;
      17'b00000000000000100: n112_o = tx_data_in;
      17'b00000000000000010: n112_o = n53_o;
      17'b00000000000000001: n112_o = tx_data_in;
      default: n112_o = tx_data_in;
    endcase
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:173:13  */
  always @*
    case (n93_o)
      17'b10000000000000000: n115_o = tx_available;
      17'b01000000000000000: n115_o = tx_available;
      17'b00100000000000000: n115_o = tx_available;
      17'b00010000000000000: n115_o = tx_available;
      17'b00001000000000000: n115_o = tx_available;
      17'b00000100000000000: n115_o = tx_available;
      17'b00000010000000000: n115_o = tx_available;
      17'b00000001000000000: n115_o = tx_available;
      17'b00000000100000000: n115_o = tx_available;
      17'b00000000010000000: n115_o = tx_available;
      17'b00000000001000000: n115_o = tx_available;
      17'b00000000000100000: n115_o = tx_available;
      17'b00000000000010000: n115_o = tx_available;
      17'b00000000000001000: n115_o = tx_available;
      17'b00000000000000100: n115_o = tx_available;
      17'b00000000000000010: n115_o = 1'b0;
      17'b00000000000000001: n115_o = 1'b1;
      default: n115_o = tx_available;
    endcase
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:173:13  */
  always @*
    case (n93_o)
      17'b10000000000000000: n133_o = 5'b00000;
      17'b01000000000000000: n133_o = 5'b10000;
      17'b00100000000000000: n133_o = 5'b01111;
      17'b00010000000000000: n133_o = 5'b01110;
      17'b00001000000000000: n133_o = 5'b01101;
      17'b00000100000000000: n133_o = 5'b01100;
      17'b00000010000000000: n133_o = 5'b01011;
      17'b00000001000000000: n133_o = 5'b01010;
      17'b00000000100000000: n133_o = 5'b01001;
      17'b00000000010000000: n133_o = 5'b01000;
      17'b00000000001000000: n133_o = 5'b00111;
      17'b00000000000100000: n133_o = 5'b00110;
      17'b00000000000010000: n133_o = 5'b00101;
      17'b00000000000001000: n133_o = 5'b00100;
      17'b00000000000000100: n133_o = 5'b00011;
      17'b00000000000000010: n133_o = 5'b00010;
      17'b00000000000000001: n133_o = n50_o;
      default: n133_o = 5'b00000;
    endcase
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:251:22  */
  assign n146_o = ~reset_btn;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:260:21  */
  assign n149_o = rdy ? 1'b1 : 1'b0;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:258:17  */
  assign n152_o = shift_state == 1'b0;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:270:17  */
  assign n154_o = shift_state == 1'b1;
  assign n155_o = {n154_o, n152_o};
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:257:13  */
  always @*
    case (n155_o)
      2'b10: n159_o = 1'b1;
      2'b01: n159_o = 1'b0;
      default: n159_o = 1'bX;
    endcase
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:257:13  */
  always @*
    case (n155_o)
      2'b10: n162_o = 1'b0;
      2'b01: n162_o = n149_o;
      default: n162_o = 1'bX;
    endcase
  assign n163_o = received_word[6:0];
  assign n164_o = output_data[6:0];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:257:13  */
  always @*
    case (n155_o)
      2'b10: n166_o = n163_o;
      2'b01: n166_o = n164_o;
      default: n166_o = 7'bX;
    endcase
  assign n167_o = received_word[7];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:257:13  */
  always @*
    case (n155_o)
      2'b10: n169_o = n167_o;
      2'b01: n169_o = 1'b0;
      default: n169_o = 1'bX;
    endcase
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:251:9  */
  assign n171_o = n146_o ? 1'b0 : n159_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:251:9  */
  assign n174_o = n146_o ? 1'b0 : 1'b1;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:251:9  */
  assign n176_o = n146_o ? 1'b0 : n162_o;
  assign n177_o = {n169_o, n166_o};
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:251:9  */
  assign n178_o = n146_o ? output_data : n177_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:280:30  */
  assign n184_o = output_data[7];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:281:30  */
  assign n185_o = output_data[6];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:282:30  */
  assign n186_o = output_data[2:0];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:297:18  */
  assign uut1_n189 = uut1_output ; // (signal)
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:294:1  */
  ros_selection uut1 (
    .challenge(mux_1_challenge),
    .enable(enable_1),
    .\output (uut1_output ));
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:305:18  */
  assign uut2_n192 = uut2_output ; // (signal)
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:302:1  */
  ros_selection uut2 (
    .challenge(mux_2_challenge),
    .enable(enable_2),
    .\output (uut2_output ));
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:312:17  */
  assign rom_n195 = rom_data_out; // (signal)
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:309:1  */
  random_rom rom (
    .address(rom_address),
    .data_out(rom_data_out));
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:332:26  */
  assign n201_o = counter_timer == 3'b001;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:334:26  */
  assign n203_o = counter_timer == 3'b010;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:336:26  */
  assign n205_o = counter_timer == 3'b011;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:338:26  */
  assign n207_o = counter_timer == 3'b100;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:338:5  */
  assign n210_o = n207_o ? 32'b00000000000000000010111011100000 : 32'b00000000000000000000000000000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:336:5  */
  assign n212_o = n205_o ? 32'b00000000000000011101010011000000 : n210_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:334:5  */
  assign n214_o = n203_o ? 32'b00000000000100100100111110000000 : n212_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:332:5  */
  assign n216_o = n201_o ? 32'b00000000101101110001101100000000 : n214_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:356:48  */
  assign n223_o = compteur_cycles + 29'b00000000000000000000000000001;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:355:9  */
  assign n225_o = enable_counter ? n223_o : 29'b00000000000000000000000000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:380:24  */
  assign n231_o = ~mode_select;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:384:45  */
  assign n232_o = rom_data_out[15:8];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:385:45  */
  assign n233_o = rom_data_out[7:0];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:380:9  */
  assign n234_o = n231_o ? internal_challenge_mux : n232_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:380:9  */
  assign n235_o = n231_o ? internal_challenge_mux : n233_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:406:36  */
  assign n236_o = ~mode_select;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:407:25  */
  assign n242_o = n496_data ? 3'b001 : 3'b100;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:413:25  */
  assign n247_o = n495_data ? 3'b001 : 3'b100;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:406:21  */
  assign n248_o = n236_o ? n242_o : n247_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:405:17  */
  assign n250_o = puf_start ? n248_o : 3'b000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:389:13  */
  assign n252_o = state == 3'b000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:433:32  */
  assign n253_o = ~mode_select;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:62  */
  assign n262_o = rom_data_out[15:8];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:62  */
  assign n267_o = rom_data_out[7:0];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:433:17  */
  assign n272_o = n253_o ? n1533_o : n3607_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:433:17  */
  assign n273_o = n253_o ? n2570_o : n4644_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:442:36  */
  assign n274_o = timer_size[30:0];  // trunc
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:442:36  */
  assign n275_o = n274_o[28:0];  // trunc
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:442:36  */
  assign n276_o = compteur_cycles == n275_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:442:17  */
  assign n279_o = n276_o ? 3'b010 : 3'b001;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:424:13  */
  assign n281_o = state == 3'b001;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:460:17  */
  assign n284_o = tx_available ? 3'b011 : 3'b010;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:448:13  */
  assign n286_o = state == 3'b010;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:475:32  */
  assign n287_o = ~mode_select;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:476:47  */
  assign n289_o = internal_challenge_mux == 8'b11111111;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:476:21  */
  assign n292_o = n289_o ? 3'b000 : 3'b100;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:482:36  */
  assign n293_o = {24'b0, rom_address};  //  uext
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:482:36  */
  assign n295_o = n293_o == 32'b00000000000000000000000011111111;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:482:21  */
  assign n298_o = n295_o ? 3'b000 : 3'b100;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:475:17  */
  assign n299_o = n287_o ? n292_o : n298_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:466:13  */
  assign n301_o = state == 3'b011;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:490:48  */
  assign n302_o = ~mode_select;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:491:90  */
  assign n304_o = internal_challenge_mux + 8'b00000001;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:493:68  */
  assign n305_o = {24'b0, rom_address};  //  uext
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:493:68  */
  assign n307_o = n305_o + 32'b00000000000000000000000000000001;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:493:56  */
  assign n308_o = n307_o[7:0];  // trunc
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:490:33  */
  assign n309_o = n302_o ? n304_o : internal_challenge_mux;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:490:33  */
  assign n310_o = n302_o ? rom_address : n308_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:489:25  */
  assign n312_o = state == 3'b100;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:508:32  */
  assign n313_o = ~mode_select;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:512:51  */
  assign n318_o = internal_challenge_mux == 8'b11111111;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:512:25  */
  assign n321_o = n318_o ? 3'b000 : 3'b100;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:509:21  */
  assign n323_o = n494_data ? 3'b001 : n321_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:522:40  */
  assign n326_o = {24'b0, rom_address};  //  uext
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:522:40  */
  assign n328_o = n326_o == 32'b00000000000000000000000011111111;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:522:25  */
  assign n331_o = n328_o ? 3'b000 : 3'b100;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:519:21  */
  assign n333_o = n493_data ? 3'b001 : n331_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:508:17  */
  assign n334_o = n313_o ? n323_o : n333_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:499:13  */
  assign n336_o = state == 3'b101;
  assign n337_o = {n336_o, n312_o, n301_o, n286_o, n281_o, n252_o};
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:388:9  */
  always @*
    case (n337_o)
      6'b100000: n344_o = 1'b0;
      6'b010000: n344_o = n489_q;
      6'b001000: n344_o = 1'b0;
      6'b000100: n344_o = 1'b1;
      6'b000010: n344_o = 1'b1;
      6'b000001: n344_o = 1'b1;
      default: n344_o = 1'bX;
    endcase
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:388:9  */
  always @*
    case (n337_o)
      6'b100000: n351_o = 1'b1;
      6'b010000: n351_o = n490_q;
      6'b001000: n351_o = 1'b0;
      6'b000100: n351_o = 1'b0;
      6'b000010: n351_o = 1'b0;
      6'b000001: n351_o = 1'b1;
      default: n351_o = 1'bX;
    endcase
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:388:9  */
  always @*
    case (n337_o)
      6'b100000: n358_o = 1'b0;
      6'b010000: n358_o = n491_q;
      6'b001000: n358_o = 1'b1;
      6'b000100: n358_o = 1'b1;
      6'b000010: n358_o = 1'b0;
      6'b000001: n358_o = 1'b1;
      default: n358_o = 1'bX;
    endcase
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:388:9  */
  always @*
    case (n337_o)
      6'b100000: n361_o = internal_challenge_mux;
      6'b010000: n361_o = n309_o;
      6'b001000: n361_o = internal_challenge_mux;
      6'b000100: n361_o = internal_challenge_mux;
      6'b000010: n361_o = internal_challenge_mux;
      6'b000001: n361_o = 8'b00000000;
      default: n361_o = 8'bX;
    endcase
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:388:9  */
  always @*
    case (n337_o)
      6'b100000: n365_o = enable_1;
      6'b010000: n365_o = enable_1;
      6'b001000: n365_o = enable_1;
      6'b000100: n365_o = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      6'b000010: n365_o = n272_o;
      6'b000001: n365_o = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      default: n365_o = 256'bX;
    endcase
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:388:9  */
  always @*
    case (n337_o)
      6'b100000: n369_o = enable_2;
      6'b010000: n369_o = enable_2;
      6'b001000: n369_o = enable_2;
      6'b000100: n369_o = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      6'b000010: n369_o = n273_o;
      6'b000001: n369_o = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      default: n369_o = 256'bX;
    endcase
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:388:9  */
  always @*
    case (n337_o)
      6'b100000: n376_o = 1'b1;
      6'b010000: n376_o = reset_counter;
      6'b001000: n376_o = 1'b0;
      6'b000100: n376_o = 1'b0;
      6'b000010: n376_o = 1'b0;
      6'b000001: n376_o = 1'b1;
      default: n376_o = 1'bX;
    endcase
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:388:9  */
  always @*
    case (n337_o)
      6'b100000: n383_o = 1'b0;
      6'b010000: n383_o = enable_comparison;
      6'b001000: n383_o = 1'b1;
      6'b000100: n383_o = 1'b0;
      6'b000010: n383_o = 1'b0;
      6'b000001: n383_o = 1'b0;
      default: n383_o = 1'bX;
    endcase
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:388:9  */
  always @*
    case (n337_o)
      6'b100000: n390_o = 1'b0;
      6'b010000: n390_o = enable_counter;
      6'b001000: n390_o = 1'b0;
      6'b000100: n390_o = 1'b0;
      6'b000010: n390_o = 1'b1;
      6'b000001: n390_o = 1'b0;
      default: n390_o = 1'bX;
    endcase
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:388:9  */
  always @*
    case (n337_o)
      6'b100000: n393_o = rom_address;
      6'b010000: n393_o = n310_o;
      6'b001000: n393_o = rom_address;
      6'b000100: n393_o = rom_address;
      6'b000010: n393_o = rom_address;
      6'b000001: n393_o = 8'b00000000;
      default: n393_o = 8'bX;
    endcase
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:388:9  */
  always @*
    case (n337_o)
      6'b100000: n396_o = n334_o;
      6'b010000: n396_o = 3'b101;
      6'b001000: n396_o = n299_o;
      6'b000100: n396_o = n284_o;
      6'b000010: n396_o = n279_o;
      6'b000001: n396_o = n250_o;
      default: n396_o = 3'bX;
    endcase
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:553:40  */
  assign n415_o = mux_2_counter + 31'b0000000000000000000000000000001;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:561:40  */
  assign n422_o = mux_1_counter + 31'b0000000000000000000000000000001;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:587:30  */
  assign n431_o = $unsigned(mux_1_counter) < $unsigned(mux_2_counter);
  assign n434_o = {mux_1_counter, mux_2_counter};
  assign n435_o = {mux_1_counter, mux_2_counter};
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:587:13  */
  assign n436_o = n431_o ? n435_o : n434_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:587:13  */
  assign n437_o = n431_o ? 1'b0 : 1'b1;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:586:9  */
  assign n444_o = enable_comparison ? 1'b1 : 1'b0;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:171:5  */
  assign n451_o = n47_o ? n111_o : tx_en;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:171:5  */
  always @(posedge clk)
    n452_q <= n451_o;
  initial
    n452_q = 1'b0;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:171:5  */
  assign n453_o = n47_o ? n112_o : tx_data_in;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:171:5  */
  always @(posedge clk)
    n454_q <= n453_o;
  initial
    n454_q = 8'b00000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:250:5  */
  always @(posedge clk)
    n455_q <= n176_o;
  initial
    n455_q = 1'b0;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:250:5  */
  always @(posedge clk)
    n456_q <= n178_o;
  initial
    n456_q = 8'b00000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:378:5  */
  always @(posedge clk)
    n457_q <= n361_o;
  initial
    n457_q = 8'b00000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:378:5  */
  assign n458_o = n18_o[63];
  assign n459_o = puf_response[63];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:585:5  */
  assign n460_o = enable_comparison ? n437_o : n459_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:585:5  */
  always @(posedge clk)
    n461_q <= n460_o;
  initial
    n461_q = n458_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:585:5  */
  assign n462_o = n18_o[61:0];
  assign n463_o = puf_response[61:0];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:585:5  */
  assign n464_o = enable_comparison ? n436_o : n463_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:585:5  */
  always @(posedge clk)
    n465_q <= n464_o;
  initial
    n465_q = n462_o;
  assign n467_o = {n461_q, 1'bZ, n465_q};
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:378:5  */
  always @(posedge clk)
    n468_q <= n234_o;
  initial
    n468_q = 8'b00000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:378:5  */
  always @(posedge clk)
    n469_q <= n235_o;
  initial
    n469_q = 8'b00000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:354:5  */
  always @(posedge clk)
    n470_q <= n225_o;
  initial
    n470_q = 29'b00000000000000000000000000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:559:1  */
  assign n471_o = enable_counter ? n422_o : mux_1_counter;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:559:1  */
  always @(posedge mux_1_out or posedge reset_counter)
    if (reset_counter)
      n472_q <= 31'b0000000000000000000000000000000;
    else
      n472_q <= n471_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:551:1  */
  assign n473_o = enable_counter ? n415_o : mux_2_counter;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:551:1  */
  always @(posedge mux_2_out or posedge reset_counter)
    if (reset_counter)
      n474_q <= 31'b0000000000000000000000000000000;
    else
      n474_q <= n473_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:378:5  */
  always @(posedge clk)
    n475_q <= n365_o;
  initial
    n475_q = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:378:5  */
  always @(posedge clk)
    n476_q <= n369_o;
  initial
    n476_q = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:378:5  */
  always @(posedge clk)
    n477_q <= n376_o;
  initial
    n477_q = 1'b0;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:378:5  */
  always @(posedge clk)
    n478_q <= n383_o;
  initial
    n478_q = 1'b0;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:378:5  */
  always @(posedge clk)
    n479_q <= n390_o;
  initial
    n479_q = 1'b0;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:585:5  */
  always @(posedge clk)
    n480_q <= n444_o;
  initial
    n480_q = 1'b1;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:171:5  */
  assign n481_o = n47_o ? n115_o : tx_available;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:171:5  */
  always @(posedge clk)
    n482_q <= n481_o;
  initial
    n482_q = 1'b1;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:378:5  */
  always @(posedge clk)
    n483_q <= n393_o;
  initial
    n483_q = 8'b00000000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:378:5  */
  always @(posedge clk)
    n484_q <= n396_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:171:5  */
  assign n485_o = n47_o ? n133_o : transmission_state;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:171:5  */
  always @(posedge clk)
    n486_q <= n485_o;
  initial
    n486_q = 5'b00000;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:250:5  */
  always @(posedge clk)
    n487_q <= n171_o;
  initial
    n487_q = 1'b0;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:250:5  */
  always @(posedge clk)
    n488_q <= n174_o;
  initial
    n488_q = 1'b0;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:378:5  */
  always @(posedge clk)
    n489_q <= n344_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:378:5  */
  always @(posedge clk)
    n490_q <= n351_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:378:5  */
  always @(posedge clk)
    n491_q <= n358_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:312:17  */
  reg n492[255:0] ; // memory
  initial begin
    n492[255] = 1'b1;
    n492[254] = 1'b1;
    n492[253] = 1'b1;
    n492[252] = 1'b1;
    n492[251] = 1'b1;
    n492[250] = 1'b1;
    n492[249] = 1'b1;
    n492[248] = 1'b1;
    n492[247] = 1'b1;
    n492[246] = 1'b1;
    n492[245] = 1'b1;
    n492[244] = 1'b1;
    n492[243] = 1'b1;
    n492[242] = 1'b1;
    n492[241] = 1'b1;
    n492[240] = 1'b1;
    n492[239] = 1'b1;
    n492[238] = 1'b1;
    n492[237] = 1'b1;
    n492[236] = 1'b1;
    n492[235] = 1'b1;
    n492[234] = 1'b1;
    n492[233] = 1'b1;
    n492[232] = 1'b1;
    n492[231] = 1'b1;
    n492[230] = 1'b1;
    n492[229] = 1'b1;
    n492[228] = 1'b1;
    n492[227] = 1'b1;
    n492[226] = 1'b1;
    n492[225] = 1'b1;
    n492[224] = 1'b1;
    n492[223] = 1'b1;
    n492[222] = 1'b1;
    n492[221] = 1'b1;
    n492[220] = 1'b1;
    n492[219] = 1'b1;
    n492[218] = 1'b1;
    n492[217] = 1'b1;
    n492[216] = 1'b1;
    n492[215] = 1'b1;
    n492[214] = 1'b1;
    n492[213] = 1'b1;
    n492[212] = 1'b1;
    n492[211] = 1'b1;
    n492[210] = 1'b1;
    n492[209] = 1'b1;
    n492[208] = 1'b1;
    n492[207] = 1'b1;
    n492[206] = 1'b1;
    n492[205] = 1'b1;
    n492[204] = 1'b1;
    n492[203] = 1'b1;
    n492[202] = 1'b1;
    n492[201] = 1'b1;
    n492[200] = 1'b1;
    n492[199] = 1'b1;
    n492[198] = 1'b1;
    n492[197] = 1'b1;
    n492[196] = 1'b1;
    n492[195] = 1'b1;
    n492[194] = 1'b1;
    n492[193] = 1'b1;
    n492[192] = 1'b1;
    n492[191] = 1'b1;
    n492[190] = 1'b1;
    n492[189] = 1'b1;
    n492[188] = 1'b1;
    n492[187] = 1'b1;
    n492[186] = 1'b1;
    n492[185] = 1'b1;
    n492[184] = 1'b1;
    n492[183] = 1'b1;
    n492[182] = 1'b1;
    n492[181] = 1'b1;
    n492[180] = 1'b1;
    n492[179] = 1'b1;
    n492[178] = 1'b1;
    n492[177] = 1'b1;
    n492[176] = 1'b1;
    n492[175] = 1'b1;
    n492[174] = 1'b1;
    n492[173] = 1'b1;
    n492[172] = 1'b1;
    n492[171] = 1'b1;
    n492[170] = 1'b1;
    n492[169] = 1'b1;
    n492[168] = 1'b1;
    n492[167] = 1'b1;
    n492[166] = 1'b1;
    n492[165] = 1'b1;
    n492[164] = 1'b1;
    n492[163] = 1'b1;
    n492[162] = 1'b1;
    n492[161] = 1'b1;
    n492[160] = 1'b1;
    n492[159] = 1'b1;
    n492[158] = 1'b1;
    n492[157] = 1'b1;
    n492[156] = 1'b1;
    n492[155] = 1'b1;
    n492[154] = 1'b1;
    n492[153] = 1'b1;
    n492[152] = 1'b1;
    n492[151] = 1'b1;
    n492[150] = 1'b1;
    n492[149] = 1'b1;
    n492[148] = 1'b1;
    n492[147] = 1'b1;
    n492[146] = 1'b1;
    n492[145] = 1'b1;
    n492[144] = 1'b1;
    n492[143] = 1'b1;
    n492[142] = 1'b1;
    n492[141] = 1'b1;
    n492[140] = 1'b1;
    n492[139] = 1'b1;
    n492[138] = 1'b1;
    n492[137] = 1'b1;
    n492[136] = 1'b1;
    n492[135] = 1'b1;
    n492[134] = 1'b1;
    n492[133] = 1'b1;
    n492[132] = 1'b1;
    n492[131] = 1'b1;
    n492[130] = 1'b1;
    n492[129] = 1'b1;
    n492[128] = 1'b1;
    n492[127] = 1'b1;
    n492[126] = 1'b1;
    n492[125] = 1'b1;
    n492[124] = 1'b1;
    n492[123] = 1'b1;
    n492[122] = 1'b1;
    n492[121] = 1'b1;
    n492[120] = 1'b1;
    n492[119] = 1'b1;
    n492[118] = 1'b1;
    n492[117] = 1'b1;
    n492[116] = 1'b1;
    n492[115] = 1'b1;
    n492[114] = 1'b1;
    n492[113] = 1'b1;
    n492[112] = 1'b1;
    n492[111] = 1'b1;
    n492[110] = 1'b1;
    n492[109] = 1'b1;
    n492[108] = 1'b1;
    n492[107] = 1'b1;
    n492[106] = 1'b1;
    n492[105] = 1'b1;
    n492[104] = 1'b1;
    n492[103] = 1'b1;
    n492[102] = 1'b1;
    n492[101] = 1'b1;
    n492[100] = 1'b1;
    n492[99] = 1'b1;
    n492[98] = 1'b1;
    n492[97] = 1'b1;
    n492[96] = 1'b1;
    n492[95] = 1'b1;
    n492[94] = 1'b1;
    n492[93] = 1'b1;
    n492[92] = 1'b1;
    n492[91] = 1'b1;
    n492[90] = 1'b1;
    n492[89] = 1'b1;
    n492[88] = 1'b1;
    n492[87] = 1'b1;
    n492[86] = 1'b1;
    n492[85] = 1'b1;
    n492[84] = 1'b1;
    n492[83] = 1'b1;
    n492[82] = 1'b1;
    n492[81] = 1'b1;
    n492[80] = 1'b1;
    n492[79] = 1'b1;
    n492[78] = 1'b1;
    n492[77] = 1'b1;
    n492[76] = 1'b1;
    n492[75] = 1'b1;
    n492[74] = 1'b1;
    n492[73] = 1'b1;
    n492[72] = 1'b1;
    n492[71] = 1'b1;
    n492[70] = 1'b1;
    n492[69] = 1'b1;
    n492[68] = 1'b1;
    n492[67] = 1'b1;
    n492[66] = 1'b1;
    n492[65] = 1'b1;
    n492[64] = 1'b1;
    n492[63] = 1'b1;
    n492[62] = 1'b1;
    n492[61] = 1'b1;
    n492[60] = 1'b1;
    n492[59] = 1'b1;
    n492[58] = 1'b1;
    n492[57] = 1'b1;
    n492[56] = 1'b1;
    n492[55] = 1'b1;
    n492[54] = 1'b1;
    n492[53] = 1'b1;
    n492[52] = 1'b1;
    n492[51] = 1'b1;
    n492[50] = 1'b1;
    n492[49] = 1'b1;
    n492[48] = 1'b1;
    n492[47] = 1'b1;
    n492[46] = 1'b1;
    n492[45] = 1'b1;
    n492[44] = 1'b1;
    n492[43] = 1'b1;
    n492[42] = 1'b1;
    n492[41] = 1'b1;
    n492[40] = 1'b1;
    n492[39] = 1'b1;
    n492[38] = 1'b1;
    n492[37] = 1'b1;
    n492[36] = 1'b1;
    n492[35] = 1'b1;
    n492[34] = 1'b1;
    n492[33] = 1'b1;
    n492[32] = 1'b1;
    n492[31] = 1'b1;
    n492[30] = 1'b1;
    n492[29] = 1'b1;
    n492[28] = 1'b1;
    n492[27] = 1'b1;
    n492[26] = 1'b1;
    n492[25] = 1'b1;
    n492[24] = 1'b1;
    n492[23] = 1'b1;
    n492[22] = 1'b1;
    n492[21] = 1'b1;
    n492[20] = 1'b1;
    n492[19] = 1'b1;
    n492[18] = 1'b1;
    n492[17] = 1'b1;
    n492[16] = 1'b1;
    n492[15] = 1'b1;
    n492[14] = 1'b1;
    n492[13] = 1'b1;
    n492[12] = 1'b1;
    n492[11] = 1'b1;
    n492[10] = 1'b1;
    n492[9] = 1'b1;
    n492[8] = 1'b1;
    n492[7] = 1'b1;
    n492[6] = 1'b1;
    n492[5] = 1'b1;
    n492[4] = 1'b1;
    n492[3] = 1'b1;
    n492[2] = 1'b1;
    n492[1] = 1'b1;
    n492[0] = 1'b1;
    end
  assign n493_data = n492[rom_address];
  assign n494_data = n492[internal_challenge_mux];
  assign n495_data = n492[rom_address];
  assign n496_data = n492[internal_challenge_mux];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:519:34  */
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:509:34  */
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:413:38  */
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:407:38  */
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n497_o = internal_challenge_mux[7];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n498_o = ~n497_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n499_o = internal_challenge_mux[6];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n500_o = ~n499_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n501_o = n498_o & n500_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n502_o = n498_o & n499_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n503_o = n497_o & n500_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n504_o = n497_o & n499_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n505_o = internal_challenge_mux[5];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n506_o = ~n505_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n507_o = n501_o & n506_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n508_o = n501_o & n505_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n509_o = n502_o & n506_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n510_o = n502_o & n505_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n511_o = n503_o & n506_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n512_o = n503_o & n505_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n513_o = n504_o & n506_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n514_o = n504_o & n505_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n515_o = internal_challenge_mux[4];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n516_o = ~n515_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n517_o = n507_o & n516_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n518_o = n507_o & n515_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n519_o = n508_o & n516_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n520_o = n508_o & n515_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n521_o = n509_o & n516_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n522_o = n509_o & n515_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n523_o = n510_o & n516_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n524_o = n510_o & n515_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n525_o = n511_o & n516_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n526_o = n511_o & n515_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n527_o = n512_o & n516_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n528_o = n512_o & n515_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n529_o = n513_o & n516_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n530_o = n513_o & n515_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n531_o = n514_o & n516_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n532_o = n514_o & n515_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n533_o = internal_challenge_mux[3];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n534_o = ~n533_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n535_o = n517_o & n534_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n536_o = n517_o & n533_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n537_o = n518_o & n534_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n538_o = n518_o & n533_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n539_o = n519_o & n534_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n540_o = n519_o & n533_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n541_o = n520_o & n534_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n542_o = n520_o & n533_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n543_o = n521_o & n534_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n544_o = n521_o & n533_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n545_o = n522_o & n534_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n546_o = n522_o & n533_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n547_o = n523_o & n534_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n548_o = n523_o & n533_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n549_o = n524_o & n534_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n550_o = n524_o & n533_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n551_o = n525_o & n534_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n552_o = n525_o & n533_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n553_o = n526_o & n534_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n554_o = n526_o & n533_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n555_o = n527_o & n534_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n556_o = n527_o & n533_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n557_o = n528_o & n534_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n558_o = n528_o & n533_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n559_o = n529_o & n534_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n560_o = n529_o & n533_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n561_o = n530_o & n534_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n562_o = n530_o & n533_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n563_o = n531_o & n534_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n564_o = n531_o & n533_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n565_o = n532_o & n534_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n566_o = n532_o & n533_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n567_o = internal_challenge_mux[2];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n568_o = ~n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n569_o = n535_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n570_o = n535_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n571_o = n536_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n572_o = n536_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n573_o = n537_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n574_o = n537_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n575_o = n538_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n576_o = n538_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n577_o = n539_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n578_o = n539_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n579_o = n540_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n580_o = n540_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n581_o = n541_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n582_o = n541_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n583_o = n542_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n584_o = n542_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n585_o = n543_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n586_o = n543_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n587_o = n544_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n588_o = n544_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n589_o = n545_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n590_o = n545_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n591_o = n546_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n592_o = n546_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n593_o = n547_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n594_o = n547_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n595_o = n548_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n596_o = n548_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n597_o = n549_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n598_o = n549_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n599_o = n550_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n600_o = n550_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n601_o = n551_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n602_o = n551_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n603_o = n552_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n604_o = n552_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n605_o = n553_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n606_o = n553_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n607_o = n554_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n608_o = n554_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n609_o = n555_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n610_o = n555_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n611_o = n556_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n612_o = n556_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n613_o = n557_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n614_o = n557_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n615_o = n558_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n616_o = n558_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n617_o = n559_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n618_o = n559_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n619_o = n560_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n620_o = n560_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n621_o = n561_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n622_o = n561_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n623_o = n562_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n624_o = n562_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n625_o = n563_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n626_o = n563_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n627_o = n564_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n628_o = n564_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n629_o = n565_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n630_o = n565_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n631_o = n566_o & n568_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n632_o = n566_o & n567_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n633_o = internal_challenge_mux[1];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n634_o = ~n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n635_o = n569_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n636_o = n569_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n637_o = n570_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n638_o = n570_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n639_o = n571_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n640_o = n571_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n641_o = n572_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n642_o = n572_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n643_o = n573_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n644_o = n573_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n645_o = n574_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n646_o = n574_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n647_o = n575_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n648_o = n575_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n649_o = n576_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n650_o = n576_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n651_o = n577_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n652_o = n577_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n653_o = n578_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n654_o = n578_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n655_o = n579_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n656_o = n579_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n657_o = n580_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n658_o = n580_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n659_o = n581_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n660_o = n581_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n661_o = n582_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n662_o = n582_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n663_o = n583_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n664_o = n583_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n665_o = n584_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n666_o = n584_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n667_o = n585_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n668_o = n585_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n669_o = n586_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n670_o = n586_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n671_o = n587_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n672_o = n587_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n673_o = n588_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n674_o = n588_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n675_o = n589_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n676_o = n589_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n677_o = n590_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n678_o = n590_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n679_o = n591_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n680_o = n591_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n681_o = n592_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n682_o = n592_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n683_o = n593_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n684_o = n593_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n685_o = n594_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n686_o = n594_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n687_o = n595_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n688_o = n595_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n689_o = n596_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n690_o = n596_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n691_o = n597_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n692_o = n597_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n693_o = n598_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n694_o = n598_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n695_o = n599_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n696_o = n599_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n697_o = n600_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n698_o = n600_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n699_o = n601_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n700_o = n601_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n701_o = n602_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n702_o = n602_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n703_o = n603_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n704_o = n603_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n705_o = n604_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n706_o = n604_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n707_o = n605_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n708_o = n605_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n709_o = n606_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n710_o = n606_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n711_o = n607_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n712_o = n607_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n713_o = n608_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n714_o = n608_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n715_o = n609_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n716_o = n609_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n717_o = n610_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n718_o = n610_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n719_o = n611_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n720_o = n611_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n721_o = n612_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n722_o = n612_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n723_o = n613_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n724_o = n613_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n725_o = n614_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n726_o = n614_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n727_o = n615_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n728_o = n615_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n729_o = n616_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n730_o = n616_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n731_o = n617_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n732_o = n617_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n733_o = n618_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n734_o = n618_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n735_o = n619_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n736_o = n619_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n737_o = n620_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n738_o = n620_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n739_o = n621_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n740_o = n621_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n741_o = n622_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n742_o = n622_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n743_o = n623_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n744_o = n623_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n745_o = n624_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n746_o = n624_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n747_o = n625_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n748_o = n625_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n749_o = n626_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n750_o = n626_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n751_o = n627_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n752_o = n627_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n753_o = n628_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n754_o = n628_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n755_o = n629_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n756_o = n629_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n757_o = n630_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n758_o = n630_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n759_o = n631_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n760_o = n631_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n761_o = n632_o & n634_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n762_o = n632_o & n633_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n763_o = internal_challenge_mux[0];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n764_o = ~n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n765_o = n635_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n766_o = n635_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n767_o = n636_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n768_o = n636_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n769_o = n637_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n770_o = n637_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n771_o = n638_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n772_o = n638_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n773_o = n639_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n774_o = n639_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n775_o = n640_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n776_o = n640_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n777_o = n641_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n778_o = n641_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n779_o = n642_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n780_o = n642_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n781_o = n643_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n782_o = n643_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n783_o = n644_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n784_o = n644_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n785_o = n645_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n786_o = n645_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n787_o = n646_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n788_o = n646_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n789_o = n647_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n790_o = n647_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n791_o = n648_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n792_o = n648_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n793_o = n649_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n794_o = n649_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n795_o = n650_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n796_o = n650_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n797_o = n651_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n798_o = n651_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n799_o = n652_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n800_o = n652_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n801_o = n653_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n802_o = n653_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n803_o = n654_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n804_o = n654_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n805_o = n655_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n806_o = n655_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n807_o = n656_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n808_o = n656_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n809_o = n657_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n810_o = n657_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n811_o = n658_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n812_o = n658_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n813_o = n659_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n814_o = n659_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n815_o = n660_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n816_o = n660_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n817_o = n661_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n818_o = n661_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n819_o = n662_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n820_o = n662_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n821_o = n663_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n822_o = n663_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n823_o = n664_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n824_o = n664_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n825_o = n665_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n826_o = n665_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n827_o = n666_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n828_o = n666_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n829_o = n667_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n830_o = n667_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n831_o = n668_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n832_o = n668_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n833_o = n669_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n834_o = n669_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n835_o = n670_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n836_o = n670_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n837_o = n671_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n838_o = n671_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n839_o = n672_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n840_o = n672_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n841_o = n673_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n842_o = n673_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n843_o = n674_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n844_o = n674_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n845_o = n675_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n846_o = n675_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n847_o = n676_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n848_o = n676_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n849_o = n677_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n850_o = n677_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n851_o = n678_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n852_o = n678_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n853_o = n679_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n854_o = n679_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n855_o = n680_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n856_o = n680_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n857_o = n681_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n858_o = n681_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n859_o = n682_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n860_o = n682_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n861_o = n683_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n862_o = n683_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n863_o = n684_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n864_o = n684_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n865_o = n685_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n866_o = n685_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n867_o = n686_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n868_o = n686_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n869_o = n687_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n870_o = n687_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n871_o = n688_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n872_o = n688_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n873_o = n689_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n874_o = n689_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n875_o = n690_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n876_o = n690_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n877_o = n691_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n878_o = n691_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n879_o = n692_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n880_o = n692_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n881_o = n693_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n882_o = n693_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n883_o = n694_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n884_o = n694_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n885_o = n695_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n886_o = n695_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n887_o = n696_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n888_o = n696_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n889_o = n697_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n890_o = n697_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n891_o = n698_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n892_o = n698_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n893_o = n699_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n894_o = n699_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n895_o = n700_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n896_o = n700_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n897_o = n701_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n898_o = n701_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n899_o = n702_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n900_o = n702_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n901_o = n703_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n902_o = n703_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n903_o = n704_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n904_o = n704_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n905_o = n705_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n906_o = n705_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n907_o = n706_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n908_o = n706_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n909_o = n707_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n910_o = n707_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n911_o = n708_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n912_o = n708_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n913_o = n709_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n914_o = n709_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n915_o = n710_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n916_o = n710_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n917_o = n711_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n918_o = n711_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n919_o = n712_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n920_o = n712_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n921_o = n713_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n922_o = n713_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n923_o = n714_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n924_o = n714_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n925_o = n715_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n926_o = n715_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n927_o = n716_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n928_o = n716_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n929_o = n717_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n930_o = n717_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n931_o = n718_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n932_o = n718_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n933_o = n719_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n934_o = n719_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n935_o = n720_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n936_o = n720_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n937_o = n721_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n938_o = n721_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n939_o = n722_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n940_o = n722_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n941_o = n723_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n942_o = n723_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n943_o = n724_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n944_o = n724_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n945_o = n725_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n946_o = n725_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n947_o = n726_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n948_o = n726_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n949_o = n727_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n950_o = n727_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n951_o = n728_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n952_o = n728_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n953_o = n729_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n954_o = n729_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n955_o = n730_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n956_o = n730_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n957_o = n731_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n958_o = n731_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n959_o = n732_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n960_o = n732_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n961_o = n733_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n962_o = n733_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n963_o = n734_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n964_o = n734_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n965_o = n735_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n966_o = n735_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n967_o = n736_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n968_o = n736_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n969_o = n737_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n970_o = n737_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n971_o = n738_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n972_o = n738_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n973_o = n739_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n974_o = n739_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n975_o = n740_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n976_o = n740_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n977_o = n741_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n978_o = n741_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n979_o = n742_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n980_o = n742_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n981_o = n743_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n982_o = n743_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n983_o = n744_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n984_o = n744_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n985_o = n745_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n986_o = n745_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n987_o = n746_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n988_o = n746_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n989_o = n747_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n990_o = n747_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n991_o = n748_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n992_o = n748_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n993_o = n749_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n994_o = n749_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n995_o = n750_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n996_o = n750_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n997_o = n751_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n998_o = n751_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n999_o = n752_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1000_o = n752_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1001_o = n753_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1002_o = n753_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1003_o = n754_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1004_o = n754_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1005_o = n755_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1006_o = n755_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1007_o = n756_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1008_o = n756_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1009_o = n757_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1010_o = n757_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1011_o = n758_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1012_o = n758_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1013_o = n759_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1014_o = n759_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1015_o = n760_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1016_o = n760_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1017_o = n761_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1018_o = n761_o & n763_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1019_o = n762_o & n764_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1020_o = n762_o & n763_o;
  assign n1021_o = enable_1[0];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1022_o = n765_o ? 1'b1 : n1021_o;
  assign n1023_o = enable_1[1];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1024_o = n766_o ? 1'b1 : n1023_o;
  assign n1025_o = enable_1[2];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1026_o = n767_o ? 1'b1 : n1025_o;
  assign n1027_o = enable_1[3];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1028_o = n768_o ? 1'b1 : n1027_o;
  assign n1029_o = enable_1[4];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1030_o = n769_o ? 1'b1 : n1029_o;
  assign n1031_o = enable_1[5];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1032_o = n770_o ? 1'b1 : n1031_o;
  assign n1033_o = enable_1[6];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1034_o = n771_o ? 1'b1 : n1033_o;
  assign n1035_o = enable_1[7];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1036_o = n772_o ? 1'b1 : n1035_o;
  assign n1037_o = enable_1[8];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1038_o = n773_o ? 1'b1 : n1037_o;
  assign n1039_o = enable_1[9];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1040_o = n774_o ? 1'b1 : n1039_o;
  assign n1041_o = enable_1[10];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1042_o = n775_o ? 1'b1 : n1041_o;
  assign n1043_o = enable_1[11];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1044_o = n776_o ? 1'b1 : n1043_o;
  assign n1045_o = enable_1[12];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1046_o = n777_o ? 1'b1 : n1045_o;
  assign n1047_o = enable_1[13];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1048_o = n778_o ? 1'b1 : n1047_o;
  assign n1049_o = enable_1[14];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1050_o = n779_o ? 1'b1 : n1049_o;
  assign n1051_o = enable_1[15];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1052_o = n780_o ? 1'b1 : n1051_o;
  assign n1053_o = enable_1[16];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1054_o = n781_o ? 1'b1 : n1053_o;
  assign n1055_o = enable_1[17];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1056_o = n782_o ? 1'b1 : n1055_o;
  assign n1057_o = enable_1[18];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1058_o = n783_o ? 1'b1 : n1057_o;
  assign n1059_o = enable_1[19];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1060_o = n784_o ? 1'b1 : n1059_o;
  assign n1061_o = enable_1[20];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1062_o = n785_o ? 1'b1 : n1061_o;
  assign n1063_o = enable_1[21];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1064_o = n786_o ? 1'b1 : n1063_o;
  assign n1065_o = enable_1[22];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1066_o = n787_o ? 1'b1 : n1065_o;
  assign n1067_o = enable_1[23];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1068_o = n788_o ? 1'b1 : n1067_o;
  assign n1069_o = enable_1[24];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1070_o = n789_o ? 1'b1 : n1069_o;
  assign n1071_o = enable_1[25];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1072_o = n790_o ? 1'b1 : n1071_o;
  assign n1073_o = enable_1[26];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1074_o = n791_o ? 1'b1 : n1073_o;
  assign n1075_o = enable_1[27];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1076_o = n792_o ? 1'b1 : n1075_o;
  assign n1077_o = enable_1[28];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1078_o = n793_o ? 1'b1 : n1077_o;
  assign n1079_o = enable_1[29];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1080_o = n794_o ? 1'b1 : n1079_o;
  assign n1081_o = enable_1[30];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1082_o = n795_o ? 1'b1 : n1081_o;
  assign n1083_o = enable_1[31];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1084_o = n796_o ? 1'b1 : n1083_o;
  assign n1085_o = enable_1[32];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1086_o = n797_o ? 1'b1 : n1085_o;
  assign n1087_o = enable_1[33];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1088_o = n798_o ? 1'b1 : n1087_o;
  assign n1089_o = enable_1[34];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1090_o = n799_o ? 1'b1 : n1089_o;
  assign n1091_o = enable_1[35];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1092_o = n800_o ? 1'b1 : n1091_o;
  assign n1093_o = enable_1[36];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1094_o = n801_o ? 1'b1 : n1093_o;
  assign n1095_o = enable_1[37];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1096_o = n802_o ? 1'b1 : n1095_o;
  assign n1097_o = enable_1[38];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1098_o = n803_o ? 1'b1 : n1097_o;
  assign n1099_o = enable_1[39];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1100_o = n804_o ? 1'b1 : n1099_o;
  assign n1101_o = enable_1[40];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1102_o = n805_o ? 1'b1 : n1101_o;
  assign n1103_o = enable_1[41];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1104_o = n806_o ? 1'b1 : n1103_o;
  assign n1105_o = enable_1[42];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1106_o = n807_o ? 1'b1 : n1105_o;
  assign n1107_o = enable_1[43];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1108_o = n808_o ? 1'b1 : n1107_o;
  assign n1109_o = enable_1[44];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1110_o = n809_o ? 1'b1 : n1109_o;
  assign n1111_o = enable_1[45];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1112_o = n810_o ? 1'b1 : n1111_o;
  assign n1113_o = enable_1[46];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1114_o = n811_o ? 1'b1 : n1113_o;
  assign n1115_o = enable_1[47];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1116_o = n812_o ? 1'b1 : n1115_o;
  assign n1117_o = enable_1[48];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1118_o = n813_o ? 1'b1 : n1117_o;
  assign n1119_o = enable_1[49];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1120_o = n814_o ? 1'b1 : n1119_o;
  assign n1121_o = enable_1[50];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1122_o = n815_o ? 1'b1 : n1121_o;
  assign n1123_o = enable_1[51];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1124_o = n816_o ? 1'b1 : n1123_o;
  assign n1125_o = enable_1[52];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1126_o = n817_o ? 1'b1 : n1125_o;
  assign n1127_o = enable_1[53];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1128_o = n818_o ? 1'b1 : n1127_o;
  assign n1129_o = enable_1[54];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1130_o = n819_o ? 1'b1 : n1129_o;
  assign n1131_o = enable_1[55];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1132_o = n820_o ? 1'b1 : n1131_o;
  assign n1133_o = enable_1[56];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1134_o = n821_o ? 1'b1 : n1133_o;
  assign n1135_o = enable_1[57];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1136_o = n822_o ? 1'b1 : n1135_o;
  assign n1137_o = enable_1[58];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1138_o = n823_o ? 1'b1 : n1137_o;
  assign n1139_o = enable_1[59];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1140_o = n824_o ? 1'b1 : n1139_o;
  assign n1141_o = enable_1[60];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1142_o = n825_o ? 1'b1 : n1141_o;
  assign n1143_o = enable_1[61];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1144_o = n826_o ? 1'b1 : n1143_o;
  assign n1145_o = enable_1[62];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1146_o = n827_o ? 1'b1 : n1145_o;
  assign n1147_o = enable_1[63];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1148_o = n828_o ? 1'b1 : n1147_o;
  assign n1149_o = enable_1[64];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1150_o = n829_o ? 1'b1 : n1149_o;
  assign n1151_o = enable_1[65];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1152_o = n830_o ? 1'b1 : n1151_o;
  assign n1153_o = enable_1[66];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1154_o = n831_o ? 1'b1 : n1153_o;
  assign n1155_o = enable_1[67];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1156_o = n832_o ? 1'b1 : n1155_o;
  assign n1157_o = enable_1[68];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1158_o = n833_o ? 1'b1 : n1157_o;
  assign n1159_o = enable_1[69];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1160_o = n834_o ? 1'b1 : n1159_o;
  assign n1161_o = enable_1[70];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1162_o = n835_o ? 1'b1 : n1161_o;
  assign n1163_o = enable_1[71];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1164_o = n836_o ? 1'b1 : n1163_o;
  assign n1165_o = enable_1[72];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1166_o = n837_o ? 1'b1 : n1165_o;
  assign n1167_o = enable_1[73];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1168_o = n838_o ? 1'b1 : n1167_o;
  assign n1169_o = enable_1[74];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1170_o = n839_o ? 1'b1 : n1169_o;
  assign n1171_o = enable_1[75];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1172_o = n840_o ? 1'b1 : n1171_o;
  assign n1173_o = enable_1[76];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1174_o = n841_o ? 1'b1 : n1173_o;
  assign n1175_o = enable_1[77];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1176_o = n842_o ? 1'b1 : n1175_o;
  assign n1177_o = enable_1[78];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1178_o = n843_o ? 1'b1 : n1177_o;
  assign n1179_o = enable_1[79];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1180_o = n844_o ? 1'b1 : n1179_o;
  assign n1181_o = enable_1[80];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1182_o = n845_o ? 1'b1 : n1181_o;
  assign n1183_o = enable_1[81];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1184_o = n846_o ? 1'b1 : n1183_o;
  assign n1185_o = enable_1[82];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1186_o = n847_o ? 1'b1 : n1185_o;
  assign n1187_o = enable_1[83];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1188_o = n848_o ? 1'b1 : n1187_o;
  assign n1189_o = enable_1[84];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1190_o = n849_o ? 1'b1 : n1189_o;
  assign n1191_o = enable_1[85];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1192_o = n850_o ? 1'b1 : n1191_o;
  assign n1193_o = enable_1[86];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1194_o = n851_o ? 1'b1 : n1193_o;
  assign n1195_o = enable_1[87];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1196_o = n852_o ? 1'b1 : n1195_o;
  assign n1197_o = enable_1[88];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1198_o = n853_o ? 1'b1 : n1197_o;
  assign n1199_o = enable_1[89];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1200_o = n854_o ? 1'b1 : n1199_o;
  assign n1201_o = enable_1[90];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1202_o = n855_o ? 1'b1 : n1201_o;
  assign n1203_o = enable_1[91];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1204_o = n856_o ? 1'b1 : n1203_o;
  assign n1205_o = enable_1[92];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1206_o = n857_o ? 1'b1 : n1205_o;
  assign n1207_o = enable_1[93];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1208_o = n858_o ? 1'b1 : n1207_o;
  assign n1209_o = enable_1[94];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1210_o = n859_o ? 1'b1 : n1209_o;
  assign n1211_o = enable_1[95];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1212_o = n860_o ? 1'b1 : n1211_o;
  assign n1213_o = enable_1[96];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1214_o = n861_o ? 1'b1 : n1213_o;
  assign n1215_o = enable_1[97];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1216_o = n862_o ? 1'b1 : n1215_o;
  assign n1217_o = enable_1[98];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1218_o = n863_o ? 1'b1 : n1217_o;
  assign n1219_o = enable_1[99];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1220_o = n864_o ? 1'b1 : n1219_o;
  assign n1221_o = enable_1[100];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1222_o = n865_o ? 1'b1 : n1221_o;
  assign n1223_o = enable_1[101];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1224_o = n866_o ? 1'b1 : n1223_o;
  assign n1225_o = enable_1[102];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1226_o = n867_o ? 1'b1 : n1225_o;
  assign n1227_o = enable_1[103];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1228_o = n868_o ? 1'b1 : n1227_o;
  assign n1229_o = enable_1[104];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1230_o = n869_o ? 1'b1 : n1229_o;
  assign n1231_o = enable_1[105];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1232_o = n870_o ? 1'b1 : n1231_o;
  assign n1233_o = enable_1[106];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1234_o = n871_o ? 1'b1 : n1233_o;
  assign n1235_o = enable_1[107];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1236_o = n872_o ? 1'b1 : n1235_o;
  assign n1237_o = enable_1[108];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1238_o = n873_o ? 1'b1 : n1237_o;
  assign n1239_o = enable_1[109];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1240_o = n874_o ? 1'b1 : n1239_o;
  assign n1241_o = enable_1[110];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1242_o = n875_o ? 1'b1 : n1241_o;
  assign n1243_o = enable_1[111];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1244_o = n876_o ? 1'b1 : n1243_o;
  assign n1245_o = enable_1[112];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1246_o = n877_o ? 1'b1 : n1245_o;
  assign n1247_o = enable_1[113];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1248_o = n878_o ? 1'b1 : n1247_o;
  assign n1249_o = enable_1[114];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1250_o = n879_o ? 1'b1 : n1249_o;
  assign n1251_o = enable_1[115];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1252_o = n880_o ? 1'b1 : n1251_o;
  assign n1253_o = enable_1[116];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1254_o = n881_o ? 1'b1 : n1253_o;
  assign n1255_o = enable_1[117];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1256_o = n882_o ? 1'b1 : n1255_o;
  assign n1257_o = enable_1[118];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1258_o = n883_o ? 1'b1 : n1257_o;
  assign n1259_o = enable_1[119];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1260_o = n884_o ? 1'b1 : n1259_o;
  assign n1261_o = enable_1[120];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1262_o = n885_o ? 1'b1 : n1261_o;
  assign n1263_o = enable_1[121];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1264_o = n886_o ? 1'b1 : n1263_o;
  assign n1265_o = enable_1[122];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1266_o = n887_o ? 1'b1 : n1265_o;
  assign n1267_o = enable_1[123];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1268_o = n888_o ? 1'b1 : n1267_o;
  assign n1269_o = enable_1[124];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1270_o = n889_o ? 1'b1 : n1269_o;
  assign n1271_o = enable_1[125];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1272_o = n890_o ? 1'b1 : n1271_o;
  assign n1273_o = enable_1[126];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1274_o = n891_o ? 1'b1 : n1273_o;
  assign n1275_o = enable_1[127];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1276_o = n892_o ? 1'b1 : n1275_o;
  assign n1277_o = enable_1[128];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1278_o = n893_o ? 1'b1 : n1277_o;
  assign n1279_o = enable_1[129];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1280_o = n894_o ? 1'b1 : n1279_o;
  assign n1281_o = enable_1[130];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1282_o = n895_o ? 1'b1 : n1281_o;
  assign n1283_o = enable_1[131];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1284_o = n896_o ? 1'b1 : n1283_o;
  assign n1285_o = enable_1[132];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1286_o = n897_o ? 1'b1 : n1285_o;
  assign n1287_o = enable_1[133];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1288_o = n898_o ? 1'b1 : n1287_o;
  assign n1289_o = enable_1[134];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1290_o = n899_o ? 1'b1 : n1289_o;
  assign n1291_o = enable_1[135];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1292_o = n900_o ? 1'b1 : n1291_o;
  assign n1293_o = enable_1[136];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1294_o = n901_o ? 1'b1 : n1293_o;
  assign n1295_o = enable_1[137];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1296_o = n902_o ? 1'b1 : n1295_o;
  assign n1297_o = enable_1[138];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1298_o = n903_o ? 1'b1 : n1297_o;
  assign n1299_o = enable_1[139];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1300_o = n904_o ? 1'b1 : n1299_o;
  assign n1301_o = enable_1[140];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1302_o = n905_o ? 1'b1 : n1301_o;
  assign n1303_o = enable_1[141];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1304_o = n906_o ? 1'b1 : n1303_o;
  assign n1305_o = enable_1[142];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1306_o = n907_o ? 1'b1 : n1305_o;
  assign n1307_o = enable_1[143];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1308_o = n908_o ? 1'b1 : n1307_o;
  assign n1309_o = enable_1[144];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1310_o = n909_o ? 1'b1 : n1309_o;
  assign n1311_o = enable_1[145];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1312_o = n910_o ? 1'b1 : n1311_o;
  assign n1313_o = enable_1[146];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1314_o = n911_o ? 1'b1 : n1313_o;
  assign n1315_o = enable_1[147];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1316_o = n912_o ? 1'b1 : n1315_o;
  assign n1317_o = enable_1[148];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1318_o = n913_o ? 1'b1 : n1317_o;
  assign n1319_o = enable_1[149];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1320_o = n914_o ? 1'b1 : n1319_o;
  assign n1321_o = enable_1[150];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1322_o = n915_o ? 1'b1 : n1321_o;
  assign n1323_o = enable_1[151];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1324_o = n916_o ? 1'b1 : n1323_o;
  assign n1325_o = enable_1[152];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1326_o = n917_o ? 1'b1 : n1325_o;
  assign n1327_o = enable_1[153];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1328_o = n918_o ? 1'b1 : n1327_o;
  assign n1329_o = enable_1[154];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1330_o = n919_o ? 1'b1 : n1329_o;
  assign n1331_o = enable_1[155];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1332_o = n920_o ? 1'b1 : n1331_o;
  assign n1333_o = enable_1[156];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1334_o = n921_o ? 1'b1 : n1333_o;
  assign n1335_o = enable_1[157];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1336_o = n922_o ? 1'b1 : n1335_o;
  assign n1337_o = enable_1[158];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1338_o = n923_o ? 1'b1 : n1337_o;
  assign n1339_o = enable_1[159];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1340_o = n924_o ? 1'b1 : n1339_o;
  assign n1341_o = enable_1[160];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1342_o = n925_o ? 1'b1 : n1341_o;
  assign n1343_o = enable_1[161];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1344_o = n926_o ? 1'b1 : n1343_o;
  assign n1345_o = enable_1[162];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1346_o = n927_o ? 1'b1 : n1345_o;
  assign n1347_o = enable_1[163];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1348_o = n928_o ? 1'b1 : n1347_o;
  assign n1349_o = enable_1[164];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1350_o = n929_o ? 1'b1 : n1349_o;
  assign n1351_o = enable_1[165];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1352_o = n930_o ? 1'b1 : n1351_o;
  assign n1353_o = enable_1[166];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1354_o = n931_o ? 1'b1 : n1353_o;
  assign n1355_o = enable_1[167];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1356_o = n932_o ? 1'b1 : n1355_o;
  assign n1357_o = enable_1[168];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1358_o = n933_o ? 1'b1 : n1357_o;
  assign n1359_o = enable_1[169];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1360_o = n934_o ? 1'b1 : n1359_o;
  assign n1361_o = enable_1[170];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1362_o = n935_o ? 1'b1 : n1361_o;
  assign n1363_o = enable_1[171];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1364_o = n936_o ? 1'b1 : n1363_o;
  assign n1365_o = enable_1[172];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1366_o = n937_o ? 1'b1 : n1365_o;
  assign n1367_o = enable_1[173];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1368_o = n938_o ? 1'b1 : n1367_o;
  assign n1369_o = enable_1[174];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1370_o = n939_o ? 1'b1 : n1369_o;
  assign n1371_o = enable_1[175];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1372_o = n940_o ? 1'b1 : n1371_o;
  assign n1373_o = enable_1[176];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1374_o = n941_o ? 1'b1 : n1373_o;
  assign n1375_o = enable_1[177];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1376_o = n942_o ? 1'b1 : n1375_o;
  assign n1377_o = enable_1[178];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1378_o = n943_o ? 1'b1 : n1377_o;
  assign n1379_o = enable_1[179];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1380_o = n944_o ? 1'b1 : n1379_o;
  assign n1381_o = enable_1[180];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1382_o = n945_o ? 1'b1 : n1381_o;
  assign n1383_o = enable_1[181];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1384_o = n946_o ? 1'b1 : n1383_o;
  assign n1385_o = enable_1[182];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1386_o = n947_o ? 1'b1 : n1385_o;
  assign n1387_o = enable_1[183];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1388_o = n948_o ? 1'b1 : n1387_o;
  assign n1389_o = enable_1[184];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1390_o = n949_o ? 1'b1 : n1389_o;
  assign n1391_o = enable_1[185];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1392_o = n950_o ? 1'b1 : n1391_o;
  assign n1393_o = enable_1[186];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1394_o = n951_o ? 1'b1 : n1393_o;
  assign n1395_o = enable_1[187];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1396_o = n952_o ? 1'b1 : n1395_o;
  assign n1397_o = enable_1[188];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1398_o = n953_o ? 1'b1 : n1397_o;
  assign n1399_o = enable_1[189];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1400_o = n954_o ? 1'b1 : n1399_o;
  assign n1401_o = enable_1[190];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1402_o = n955_o ? 1'b1 : n1401_o;
  assign n1403_o = enable_1[191];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1404_o = n956_o ? 1'b1 : n1403_o;
  assign n1405_o = enable_1[192];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1406_o = n957_o ? 1'b1 : n1405_o;
  assign n1407_o = enable_1[193];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1408_o = n958_o ? 1'b1 : n1407_o;
  assign n1409_o = enable_1[194];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1410_o = n959_o ? 1'b1 : n1409_o;
  assign n1411_o = enable_1[195];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1412_o = n960_o ? 1'b1 : n1411_o;
  assign n1413_o = enable_1[196];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1414_o = n961_o ? 1'b1 : n1413_o;
  assign n1415_o = enable_1[197];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1416_o = n962_o ? 1'b1 : n1415_o;
  assign n1417_o = enable_1[198];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1418_o = n963_o ? 1'b1 : n1417_o;
  assign n1419_o = enable_1[199];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1420_o = n964_o ? 1'b1 : n1419_o;
  assign n1421_o = enable_1[200];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1422_o = n965_o ? 1'b1 : n1421_o;
  assign n1423_o = enable_1[201];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1424_o = n966_o ? 1'b1 : n1423_o;
  assign n1425_o = enable_1[202];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1426_o = n967_o ? 1'b1 : n1425_o;
  assign n1427_o = enable_1[203];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1428_o = n968_o ? 1'b1 : n1427_o;
  assign n1429_o = enable_1[204];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1430_o = n969_o ? 1'b1 : n1429_o;
  assign n1431_o = enable_1[205];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1432_o = n970_o ? 1'b1 : n1431_o;
  assign n1433_o = enable_1[206];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1434_o = n971_o ? 1'b1 : n1433_o;
  assign n1435_o = enable_1[207];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1436_o = n972_o ? 1'b1 : n1435_o;
  assign n1437_o = enable_1[208];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1438_o = n973_o ? 1'b1 : n1437_o;
  assign n1439_o = enable_1[209];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1440_o = n974_o ? 1'b1 : n1439_o;
  assign n1441_o = enable_1[210];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1442_o = n975_o ? 1'b1 : n1441_o;
  assign n1443_o = enable_1[211];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1444_o = n976_o ? 1'b1 : n1443_o;
  assign n1445_o = enable_1[212];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1446_o = n977_o ? 1'b1 : n1445_o;
  assign n1447_o = enable_1[213];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1448_o = n978_o ? 1'b1 : n1447_o;
  assign n1449_o = enable_1[214];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1450_o = n979_o ? 1'b1 : n1449_o;
  assign n1451_o = enable_1[215];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1452_o = n980_o ? 1'b1 : n1451_o;
  assign n1453_o = enable_1[216];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1454_o = n981_o ? 1'b1 : n1453_o;
  assign n1455_o = enable_1[217];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1456_o = n982_o ? 1'b1 : n1455_o;
  assign n1457_o = enable_1[218];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1458_o = n983_o ? 1'b1 : n1457_o;
  assign n1459_o = enable_1[219];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1460_o = n984_o ? 1'b1 : n1459_o;
  assign n1461_o = enable_1[220];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1462_o = n985_o ? 1'b1 : n1461_o;
  assign n1463_o = enable_1[221];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1464_o = n986_o ? 1'b1 : n1463_o;
  assign n1465_o = enable_1[222];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1466_o = n987_o ? 1'b1 : n1465_o;
  assign n1467_o = enable_1[223];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1468_o = n988_o ? 1'b1 : n1467_o;
  assign n1469_o = enable_1[224];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1470_o = n989_o ? 1'b1 : n1469_o;
  assign n1471_o = enable_1[225];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1472_o = n990_o ? 1'b1 : n1471_o;
  assign n1473_o = enable_1[226];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1474_o = n991_o ? 1'b1 : n1473_o;
  assign n1475_o = enable_1[227];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1476_o = n992_o ? 1'b1 : n1475_o;
  assign n1477_o = enable_1[228];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1478_o = n993_o ? 1'b1 : n1477_o;
  assign n1479_o = enable_1[229];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1480_o = n994_o ? 1'b1 : n1479_o;
  assign n1481_o = enable_1[230];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1482_o = n995_o ? 1'b1 : n1481_o;
  assign n1483_o = enable_1[231];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1484_o = n996_o ? 1'b1 : n1483_o;
  assign n1485_o = enable_1[232];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1486_o = n997_o ? 1'b1 : n1485_o;
  assign n1487_o = enable_1[233];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1488_o = n998_o ? 1'b1 : n1487_o;
  assign n1489_o = enable_1[234];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1490_o = n999_o ? 1'b1 : n1489_o;
  assign n1491_o = enable_1[235];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1492_o = n1000_o ? 1'b1 : n1491_o;
  assign n1493_o = enable_1[236];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1494_o = n1001_o ? 1'b1 : n1493_o;
  assign n1495_o = enable_1[237];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1496_o = n1002_o ? 1'b1 : n1495_o;
  assign n1497_o = enable_1[238];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1498_o = n1003_o ? 1'b1 : n1497_o;
  assign n1499_o = enable_1[239];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1500_o = n1004_o ? 1'b1 : n1499_o;
  assign n1501_o = enable_1[240];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1502_o = n1005_o ? 1'b1 : n1501_o;
  assign n1503_o = enable_1[241];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1504_o = n1006_o ? 1'b1 : n1503_o;
  assign n1505_o = enable_1[242];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1506_o = n1007_o ? 1'b1 : n1505_o;
  assign n1507_o = enable_1[243];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1508_o = n1008_o ? 1'b1 : n1507_o;
  assign n1509_o = enable_1[244];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1510_o = n1009_o ? 1'b1 : n1509_o;
  assign n1511_o = enable_1[245];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1512_o = n1010_o ? 1'b1 : n1511_o;
  assign n1513_o = enable_1[246];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1514_o = n1011_o ? 1'b1 : n1513_o;
  assign n1515_o = enable_1[247];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1516_o = n1012_o ? 1'b1 : n1515_o;
  assign n1517_o = enable_1[248];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1518_o = n1013_o ? 1'b1 : n1517_o;
  assign n1519_o = enable_1[249];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1520_o = n1014_o ? 1'b1 : n1519_o;
  assign n1521_o = enable_1[250];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1522_o = n1015_o ? 1'b1 : n1521_o;
  assign n1523_o = enable_1[251];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1524_o = n1016_o ? 1'b1 : n1523_o;
  assign n1525_o = enable_1[252];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1526_o = n1017_o ? 1'b1 : n1525_o;
  assign n1527_o = enable_1[253];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1528_o = n1018_o ? 1'b1 : n1527_o;
  assign n1529_o = enable_1[254];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1530_o = n1019_o ? 1'b1 : n1529_o;
  assign n1531_o = enable_1[255];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:434:21  */
  assign n1532_o = n1020_o ? 1'b1 : n1531_o;
  assign n1533_o = {n1532_o, n1530_o, n1528_o, n1526_o, n1524_o, n1522_o, n1520_o, n1518_o, n1516_o, n1514_o, n1512_o, n1510_o, n1508_o, n1506_o, n1504_o, n1502_o, n1500_o, n1498_o, n1496_o, n1494_o, n1492_o, n1490_o, n1488_o, n1486_o, n1484_o, n1482_o, n1480_o, n1478_o, n1476_o, n1474_o, n1472_o, n1470_o, n1468_o, n1466_o, n1464_o, n1462_o, n1460_o, n1458_o, n1456_o, n1454_o, n1452_o, n1450_o, n1448_o, n1446_o, n1444_o, n1442_o, n1440_o, n1438_o, n1436_o, n1434_o, n1432_o, n1430_o, n1428_o, n1426_o, n1424_o, n1422_o, n1420_o, n1418_o, n1416_o, n1414_o, n1412_o, n1410_o, n1408_o, n1406_o, n1404_o, n1402_o, n1400_o, n1398_o, n1396_o, n1394_o, n1392_o, n1390_o, n1388_o, n1386_o, n1384_o, n1382_o, n1380_o, n1378_o, n1376_o, n1374_o, n1372_o, n1370_o, n1368_o, n1366_o, n1364_o, n1362_o, n1360_o, n1358_o, n1356_o, n1354_o, n1352_o, n1350_o, n1348_o, n1346_o, n1344_o, n1342_o, n1340_o, n1338_o, n1336_o, n1334_o, n1332_o, n1330_o, n1328_o, n1326_o, n1324_o, n1322_o, n1320_o, n1318_o, n1316_o, n1314_o, n1312_o, n1310_o, n1308_o, n1306_o, n1304_o, n1302_o, n1300_o, n1298_o, n1296_o, n1294_o, n1292_o, n1290_o, n1288_o, n1286_o, n1284_o, n1282_o, n1280_o, n1278_o, n1276_o, n1274_o, n1272_o, n1270_o, n1268_o, n1266_o, n1264_o, n1262_o, n1260_o, n1258_o, n1256_o, n1254_o, n1252_o, n1250_o, n1248_o, n1246_o, n1244_o, n1242_o, n1240_o, n1238_o, n1236_o, n1234_o, n1232_o, n1230_o, n1228_o, n1226_o, n1224_o, n1222_o, n1220_o, n1218_o, n1216_o, n1214_o, n1212_o, n1210_o, n1208_o, n1206_o, n1204_o, n1202_o, n1200_o, n1198_o, n1196_o, n1194_o, n1192_o, n1190_o, n1188_o, n1186_o, n1184_o, n1182_o, n1180_o, n1178_o, n1176_o, n1174_o, n1172_o, n1170_o, n1168_o, n1166_o, n1164_o, n1162_o, n1160_o, n1158_o, n1156_o, n1154_o, n1152_o, n1150_o, n1148_o, n1146_o, n1144_o, n1142_o, n1140_o, n1138_o, n1136_o, n1134_o, n1132_o, n1130_o, n1128_o, n1126_o, n1124_o, n1122_o, n1120_o, n1118_o, n1116_o, n1114_o, n1112_o, n1110_o, n1108_o, n1106_o, n1104_o, n1102_o, n1100_o, n1098_o, n1096_o, n1094_o, n1092_o, n1090_o, n1088_o, n1086_o, n1084_o, n1082_o, n1080_o, n1078_o, n1076_o, n1074_o, n1072_o, n1070_o, n1068_o, n1066_o, n1064_o, n1062_o, n1060_o, n1058_o, n1056_o, n1054_o, n1052_o, n1050_o, n1048_o, n1046_o, n1044_o, n1042_o, n1040_o, n1038_o, n1036_o, n1034_o, n1032_o, n1030_o, n1028_o, n1026_o, n1024_o, n1022_o};
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1534_o = internal_challenge_mux[7];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1535_o = ~n1534_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1536_o = internal_challenge_mux[6];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1537_o = ~n1536_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1538_o = n1535_o & n1537_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1539_o = n1535_o & n1536_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1540_o = n1534_o & n1537_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1541_o = n1534_o & n1536_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1542_o = internal_challenge_mux[5];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1543_o = ~n1542_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1544_o = n1538_o & n1543_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1545_o = n1538_o & n1542_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1546_o = n1539_o & n1543_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1547_o = n1539_o & n1542_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1548_o = n1540_o & n1543_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1549_o = n1540_o & n1542_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1550_o = n1541_o & n1543_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1551_o = n1541_o & n1542_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1552_o = internal_challenge_mux[4];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1553_o = ~n1552_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1554_o = n1544_o & n1553_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1555_o = n1544_o & n1552_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1556_o = n1545_o & n1553_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1557_o = n1545_o & n1552_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1558_o = n1546_o & n1553_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1559_o = n1546_o & n1552_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1560_o = n1547_o & n1553_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1561_o = n1547_o & n1552_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1562_o = n1548_o & n1553_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1563_o = n1548_o & n1552_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1564_o = n1549_o & n1553_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1565_o = n1549_o & n1552_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1566_o = n1550_o & n1553_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1567_o = n1550_o & n1552_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1568_o = n1551_o & n1553_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1569_o = n1551_o & n1552_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1570_o = internal_challenge_mux[3];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1571_o = ~n1570_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1572_o = n1554_o & n1571_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1573_o = n1554_o & n1570_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1574_o = n1555_o & n1571_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1575_o = n1555_o & n1570_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1576_o = n1556_o & n1571_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1577_o = n1556_o & n1570_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1578_o = n1557_o & n1571_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1579_o = n1557_o & n1570_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1580_o = n1558_o & n1571_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1581_o = n1558_o & n1570_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1582_o = n1559_o & n1571_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1583_o = n1559_o & n1570_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1584_o = n1560_o & n1571_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1585_o = n1560_o & n1570_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1586_o = n1561_o & n1571_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1587_o = n1561_o & n1570_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1588_o = n1562_o & n1571_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1589_o = n1562_o & n1570_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1590_o = n1563_o & n1571_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1591_o = n1563_o & n1570_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1592_o = n1564_o & n1571_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1593_o = n1564_o & n1570_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1594_o = n1565_o & n1571_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1595_o = n1565_o & n1570_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1596_o = n1566_o & n1571_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1597_o = n1566_o & n1570_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1598_o = n1567_o & n1571_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1599_o = n1567_o & n1570_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1600_o = n1568_o & n1571_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1601_o = n1568_o & n1570_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1602_o = n1569_o & n1571_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1603_o = n1569_o & n1570_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1604_o = internal_challenge_mux[2];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1605_o = ~n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1606_o = n1572_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1607_o = n1572_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1608_o = n1573_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1609_o = n1573_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1610_o = n1574_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1611_o = n1574_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1612_o = n1575_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1613_o = n1575_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1614_o = n1576_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1615_o = n1576_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1616_o = n1577_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1617_o = n1577_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1618_o = n1578_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1619_o = n1578_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1620_o = n1579_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1621_o = n1579_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1622_o = n1580_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1623_o = n1580_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1624_o = n1581_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1625_o = n1581_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1626_o = n1582_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1627_o = n1582_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1628_o = n1583_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1629_o = n1583_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1630_o = n1584_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1631_o = n1584_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1632_o = n1585_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1633_o = n1585_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1634_o = n1586_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1635_o = n1586_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1636_o = n1587_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1637_o = n1587_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1638_o = n1588_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1639_o = n1588_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1640_o = n1589_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1641_o = n1589_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1642_o = n1590_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1643_o = n1590_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1644_o = n1591_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1645_o = n1591_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1646_o = n1592_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1647_o = n1592_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1648_o = n1593_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1649_o = n1593_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1650_o = n1594_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1651_o = n1594_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1652_o = n1595_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1653_o = n1595_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1654_o = n1596_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1655_o = n1596_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1656_o = n1597_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1657_o = n1597_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1658_o = n1598_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1659_o = n1598_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1660_o = n1599_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1661_o = n1599_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1662_o = n1600_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1663_o = n1600_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1664_o = n1601_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1665_o = n1601_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1666_o = n1602_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1667_o = n1602_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1668_o = n1603_o & n1605_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1669_o = n1603_o & n1604_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1670_o = internal_challenge_mux[1];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1671_o = ~n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1672_o = n1606_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1673_o = n1606_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1674_o = n1607_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1675_o = n1607_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1676_o = n1608_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1677_o = n1608_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1678_o = n1609_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1679_o = n1609_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1680_o = n1610_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1681_o = n1610_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1682_o = n1611_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1683_o = n1611_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1684_o = n1612_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1685_o = n1612_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1686_o = n1613_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1687_o = n1613_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1688_o = n1614_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1689_o = n1614_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1690_o = n1615_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1691_o = n1615_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1692_o = n1616_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1693_o = n1616_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1694_o = n1617_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1695_o = n1617_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1696_o = n1618_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1697_o = n1618_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1698_o = n1619_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1699_o = n1619_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1700_o = n1620_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1701_o = n1620_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1702_o = n1621_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1703_o = n1621_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1704_o = n1622_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1705_o = n1622_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1706_o = n1623_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1707_o = n1623_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1708_o = n1624_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1709_o = n1624_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1710_o = n1625_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1711_o = n1625_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1712_o = n1626_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1713_o = n1626_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1714_o = n1627_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1715_o = n1627_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1716_o = n1628_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1717_o = n1628_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1718_o = n1629_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1719_o = n1629_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1720_o = n1630_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1721_o = n1630_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1722_o = n1631_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1723_o = n1631_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1724_o = n1632_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1725_o = n1632_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1726_o = n1633_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1727_o = n1633_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1728_o = n1634_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1729_o = n1634_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1730_o = n1635_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1731_o = n1635_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1732_o = n1636_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1733_o = n1636_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1734_o = n1637_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1735_o = n1637_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1736_o = n1638_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1737_o = n1638_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1738_o = n1639_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1739_o = n1639_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1740_o = n1640_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1741_o = n1640_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1742_o = n1641_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1743_o = n1641_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1744_o = n1642_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1745_o = n1642_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1746_o = n1643_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1747_o = n1643_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1748_o = n1644_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1749_o = n1644_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1750_o = n1645_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1751_o = n1645_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1752_o = n1646_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1753_o = n1646_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1754_o = n1647_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1755_o = n1647_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1756_o = n1648_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1757_o = n1648_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1758_o = n1649_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1759_o = n1649_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1760_o = n1650_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1761_o = n1650_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1762_o = n1651_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1763_o = n1651_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1764_o = n1652_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1765_o = n1652_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1766_o = n1653_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1767_o = n1653_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1768_o = n1654_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1769_o = n1654_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1770_o = n1655_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1771_o = n1655_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1772_o = n1656_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1773_o = n1656_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1774_o = n1657_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1775_o = n1657_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1776_o = n1658_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1777_o = n1658_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1778_o = n1659_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1779_o = n1659_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1780_o = n1660_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1781_o = n1660_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1782_o = n1661_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1783_o = n1661_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1784_o = n1662_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1785_o = n1662_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1786_o = n1663_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1787_o = n1663_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1788_o = n1664_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1789_o = n1664_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1790_o = n1665_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1791_o = n1665_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1792_o = n1666_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1793_o = n1666_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1794_o = n1667_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1795_o = n1667_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1796_o = n1668_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1797_o = n1668_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1798_o = n1669_o & n1671_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1799_o = n1669_o & n1670_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1800_o = internal_challenge_mux[0];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1801_o = ~n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1802_o = n1672_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1803_o = n1672_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1804_o = n1673_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1805_o = n1673_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1806_o = n1674_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1807_o = n1674_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1808_o = n1675_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1809_o = n1675_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1810_o = n1676_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1811_o = n1676_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1812_o = n1677_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1813_o = n1677_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1814_o = n1678_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1815_o = n1678_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1816_o = n1679_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1817_o = n1679_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1818_o = n1680_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1819_o = n1680_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1820_o = n1681_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1821_o = n1681_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1822_o = n1682_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1823_o = n1682_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1824_o = n1683_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1825_o = n1683_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1826_o = n1684_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1827_o = n1684_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1828_o = n1685_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1829_o = n1685_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1830_o = n1686_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1831_o = n1686_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1832_o = n1687_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1833_o = n1687_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1834_o = n1688_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1835_o = n1688_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1836_o = n1689_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1837_o = n1689_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1838_o = n1690_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1839_o = n1690_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1840_o = n1691_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1841_o = n1691_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1842_o = n1692_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1843_o = n1692_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1844_o = n1693_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1845_o = n1693_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1846_o = n1694_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1847_o = n1694_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1848_o = n1695_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1849_o = n1695_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1850_o = n1696_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1851_o = n1696_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1852_o = n1697_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1853_o = n1697_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1854_o = n1698_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1855_o = n1698_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1856_o = n1699_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1857_o = n1699_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1858_o = n1700_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1859_o = n1700_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1860_o = n1701_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1861_o = n1701_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1862_o = n1702_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1863_o = n1702_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1864_o = n1703_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1865_o = n1703_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1866_o = n1704_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1867_o = n1704_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1868_o = n1705_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1869_o = n1705_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1870_o = n1706_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1871_o = n1706_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1872_o = n1707_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1873_o = n1707_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1874_o = n1708_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1875_o = n1708_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1876_o = n1709_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1877_o = n1709_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1878_o = n1710_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1879_o = n1710_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1880_o = n1711_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1881_o = n1711_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1882_o = n1712_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1883_o = n1712_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1884_o = n1713_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1885_o = n1713_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1886_o = n1714_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1887_o = n1714_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1888_o = n1715_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1889_o = n1715_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1890_o = n1716_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1891_o = n1716_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1892_o = n1717_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1893_o = n1717_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1894_o = n1718_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1895_o = n1718_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1896_o = n1719_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1897_o = n1719_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1898_o = n1720_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1899_o = n1720_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1900_o = n1721_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1901_o = n1721_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1902_o = n1722_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1903_o = n1722_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1904_o = n1723_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1905_o = n1723_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1906_o = n1724_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1907_o = n1724_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1908_o = n1725_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1909_o = n1725_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1910_o = n1726_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1911_o = n1726_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1912_o = n1727_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1913_o = n1727_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1914_o = n1728_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1915_o = n1728_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1916_o = n1729_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1917_o = n1729_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1918_o = n1730_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1919_o = n1730_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1920_o = n1731_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1921_o = n1731_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1922_o = n1732_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1923_o = n1732_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1924_o = n1733_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1925_o = n1733_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1926_o = n1734_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1927_o = n1734_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1928_o = n1735_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1929_o = n1735_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1930_o = n1736_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1931_o = n1736_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1932_o = n1737_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1933_o = n1737_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1934_o = n1738_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1935_o = n1738_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1936_o = n1739_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1937_o = n1739_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1938_o = n1740_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1939_o = n1740_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1940_o = n1741_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1941_o = n1741_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1942_o = n1742_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1943_o = n1742_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1944_o = n1743_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1945_o = n1743_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1946_o = n1744_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1947_o = n1744_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1948_o = n1745_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1949_o = n1745_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1950_o = n1746_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1951_o = n1746_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1952_o = n1747_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1953_o = n1747_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1954_o = n1748_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1955_o = n1748_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1956_o = n1749_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1957_o = n1749_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1958_o = n1750_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1959_o = n1750_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1960_o = n1751_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1961_o = n1751_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1962_o = n1752_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1963_o = n1752_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1964_o = n1753_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1965_o = n1753_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1966_o = n1754_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1967_o = n1754_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1968_o = n1755_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1969_o = n1755_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1970_o = n1756_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1971_o = n1756_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1972_o = n1757_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1973_o = n1757_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1974_o = n1758_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1975_o = n1758_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1976_o = n1759_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1977_o = n1759_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1978_o = n1760_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1979_o = n1760_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1980_o = n1761_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1981_o = n1761_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1982_o = n1762_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1983_o = n1762_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1984_o = n1763_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1985_o = n1763_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1986_o = n1764_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1987_o = n1764_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1988_o = n1765_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1989_o = n1765_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1990_o = n1766_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1991_o = n1766_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1992_o = n1767_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1993_o = n1767_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1994_o = n1768_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1995_o = n1768_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1996_o = n1769_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1997_o = n1769_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1998_o = n1770_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n1999_o = n1770_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2000_o = n1771_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2001_o = n1771_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2002_o = n1772_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2003_o = n1772_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2004_o = n1773_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2005_o = n1773_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2006_o = n1774_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2007_o = n1774_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2008_o = n1775_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2009_o = n1775_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2010_o = n1776_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2011_o = n1776_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2012_o = n1777_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2013_o = n1777_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2014_o = n1778_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2015_o = n1778_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2016_o = n1779_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2017_o = n1779_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2018_o = n1780_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2019_o = n1780_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2020_o = n1781_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2021_o = n1781_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2022_o = n1782_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2023_o = n1782_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2024_o = n1783_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2025_o = n1783_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2026_o = n1784_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2027_o = n1784_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2028_o = n1785_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2029_o = n1785_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2030_o = n1786_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2031_o = n1786_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2032_o = n1787_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2033_o = n1787_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2034_o = n1788_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2035_o = n1788_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2036_o = n1789_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2037_o = n1789_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2038_o = n1790_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2039_o = n1790_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2040_o = n1791_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2041_o = n1791_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2042_o = n1792_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2043_o = n1792_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2044_o = n1793_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2045_o = n1793_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2046_o = n1794_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2047_o = n1794_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2048_o = n1795_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2049_o = n1795_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2050_o = n1796_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2051_o = n1796_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2052_o = n1797_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2053_o = n1797_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2054_o = n1798_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2055_o = n1798_o & n1800_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2056_o = n1799_o & n1801_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2057_o = n1799_o & n1800_o;
  assign n2058_o = enable_2[0];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2059_o = n1802_o ? 1'b1 : n2058_o;
  assign n2060_o = enable_2[1];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2061_o = n1803_o ? 1'b1 : n2060_o;
  assign n2062_o = enable_2[2];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2063_o = n1804_o ? 1'b1 : n2062_o;
  assign n2064_o = enable_2[3];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2065_o = n1805_o ? 1'b1 : n2064_o;
  assign n2066_o = enable_2[4];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2067_o = n1806_o ? 1'b1 : n2066_o;
  assign n2068_o = enable_2[5];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2069_o = n1807_o ? 1'b1 : n2068_o;
  assign n2070_o = enable_2[6];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2071_o = n1808_o ? 1'b1 : n2070_o;
  assign n2072_o = enable_2[7];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2073_o = n1809_o ? 1'b1 : n2072_o;
  assign n2074_o = enable_2[8];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2075_o = n1810_o ? 1'b1 : n2074_o;
  assign n2076_o = enable_2[9];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2077_o = n1811_o ? 1'b1 : n2076_o;
  assign n2078_o = enable_2[10];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2079_o = n1812_o ? 1'b1 : n2078_o;
  assign n2080_o = enable_2[11];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2081_o = n1813_o ? 1'b1 : n2080_o;
  assign n2082_o = enable_2[12];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2083_o = n1814_o ? 1'b1 : n2082_o;
  assign n2084_o = enable_2[13];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2085_o = n1815_o ? 1'b1 : n2084_o;
  assign n2086_o = enable_2[14];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2087_o = n1816_o ? 1'b1 : n2086_o;
  assign n2088_o = enable_2[15];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2089_o = n1817_o ? 1'b1 : n2088_o;
  assign n2090_o = enable_2[16];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2091_o = n1818_o ? 1'b1 : n2090_o;
  assign n2092_o = enable_2[17];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2093_o = n1819_o ? 1'b1 : n2092_o;
  assign n2094_o = enable_2[18];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2095_o = n1820_o ? 1'b1 : n2094_o;
  assign n2096_o = enable_2[19];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2097_o = n1821_o ? 1'b1 : n2096_o;
  assign n2098_o = enable_2[20];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2099_o = n1822_o ? 1'b1 : n2098_o;
  assign n2100_o = enable_2[21];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2101_o = n1823_o ? 1'b1 : n2100_o;
  assign n2102_o = enable_2[22];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2103_o = n1824_o ? 1'b1 : n2102_o;
  assign n2104_o = enable_2[23];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2105_o = n1825_o ? 1'b1 : n2104_o;
  assign n2106_o = enable_2[24];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2107_o = n1826_o ? 1'b1 : n2106_o;
  assign n2108_o = enable_2[25];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2109_o = n1827_o ? 1'b1 : n2108_o;
  assign n2110_o = enable_2[26];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2111_o = n1828_o ? 1'b1 : n2110_o;
  assign n2112_o = enable_2[27];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2113_o = n1829_o ? 1'b1 : n2112_o;
  assign n2114_o = enable_2[28];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2115_o = n1830_o ? 1'b1 : n2114_o;
  assign n2116_o = enable_2[29];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2117_o = n1831_o ? 1'b1 : n2116_o;
  assign n2118_o = enable_2[30];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2119_o = n1832_o ? 1'b1 : n2118_o;
  assign n2120_o = enable_2[31];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2121_o = n1833_o ? 1'b1 : n2120_o;
  assign n2122_o = enable_2[32];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2123_o = n1834_o ? 1'b1 : n2122_o;
  assign n2124_o = enable_2[33];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2125_o = n1835_o ? 1'b1 : n2124_o;
  assign n2126_o = enable_2[34];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2127_o = n1836_o ? 1'b1 : n2126_o;
  assign n2128_o = enable_2[35];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2129_o = n1837_o ? 1'b1 : n2128_o;
  assign n2130_o = enable_2[36];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2131_o = n1838_o ? 1'b1 : n2130_o;
  assign n2132_o = enable_2[37];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2133_o = n1839_o ? 1'b1 : n2132_o;
  assign n2134_o = enable_2[38];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2135_o = n1840_o ? 1'b1 : n2134_o;
  assign n2136_o = enable_2[39];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2137_o = n1841_o ? 1'b1 : n2136_o;
  assign n2138_o = enable_2[40];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2139_o = n1842_o ? 1'b1 : n2138_o;
  assign n2140_o = enable_2[41];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2141_o = n1843_o ? 1'b1 : n2140_o;
  assign n2142_o = enable_2[42];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2143_o = n1844_o ? 1'b1 : n2142_o;
  assign n2144_o = enable_2[43];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2145_o = n1845_o ? 1'b1 : n2144_o;
  assign n2146_o = enable_2[44];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2147_o = n1846_o ? 1'b1 : n2146_o;
  assign n2148_o = enable_2[45];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2149_o = n1847_o ? 1'b1 : n2148_o;
  assign n2150_o = enable_2[46];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2151_o = n1848_o ? 1'b1 : n2150_o;
  assign n2152_o = enable_2[47];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2153_o = n1849_o ? 1'b1 : n2152_o;
  assign n2154_o = enable_2[48];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2155_o = n1850_o ? 1'b1 : n2154_o;
  assign n2156_o = enable_2[49];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2157_o = n1851_o ? 1'b1 : n2156_o;
  assign n2158_o = enable_2[50];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2159_o = n1852_o ? 1'b1 : n2158_o;
  assign n2160_o = enable_2[51];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2161_o = n1853_o ? 1'b1 : n2160_o;
  assign n2162_o = enable_2[52];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2163_o = n1854_o ? 1'b1 : n2162_o;
  assign n2164_o = enable_2[53];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2165_o = n1855_o ? 1'b1 : n2164_o;
  assign n2166_o = enable_2[54];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2167_o = n1856_o ? 1'b1 : n2166_o;
  assign n2168_o = enable_2[55];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2169_o = n1857_o ? 1'b1 : n2168_o;
  assign n2170_o = enable_2[56];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2171_o = n1858_o ? 1'b1 : n2170_o;
  assign n2172_o = enable_2[57];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2173_o = n1859_o ? 1'b1 : n2172_o;
  assign n2174_o = enable_2[58];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2175_o = n1860_o ? 1'b1 : n2174_o;
  assign n2176_o = enable_2[59];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2177_o = n1861_o ? 1'b1 : n2176_o;
  assign n2178_o = enable_2[60];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2179_o = n1862_o ? 1'b1 : n2178_o;
  assign n2180_o = enable_2[61];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2181_o = n1863_o ? 1'b1 : n2180_o;
  assign n2182_o = enable_2[62];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2183_o = n1864_o ? 1'b1 : n2182_o;
  assign n2184_o = enable_2[63];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2185_o = n1865_o ? 1'b1 : n2184_o;
  assign n2186_o = enable_2[64];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2187_o = n1866_o ? 1'b1 : n2186_o;
  assign n2188_o = enable_2[65];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2189_o = n1867_o ? 1'b1 : n2188_o;
  assign n2190_o = enable_2[66];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2191_o = n1868_o ? 1'b1 : n2190_o;
  assign n2192_o = enable_2[67];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2193_o = n1869_o ? 1'b1 : n2192_o;
  assign n2194_o = enable_2[68];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2195_o = n1870_o ? 1'b1 : n2194_o;
  assign n2196_o = enable_2[69];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2197_o = n1871_o ? 1'b1 : n2196_o;
  assign n2198_o = enable_2[70];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2199_o = n1872_o ? 1'b1 : n2198_o;
  assign n2200_o = enable_2[71];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2201_o = n1873_o ? 1'b1 : n2200_o;
  assign n2202_o = enable_2[72];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2203_o = n1874_o ? 1'b1 : n2202_o;
  assign n2204_o = enable_2[73];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2205_o = n1875_o ? 1'b1 : n2204_o;
  assign n2206_o = enable_2[74];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2207_o = n1876_o ? 1'b1 : n2206_o;
  assign n2208_o = enable_2[75];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2209_o = n1877_o ? 1'b1 : n2208_o;
  assign n2210_o = enable_2[76];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2211_o = n1878_o ? 1'b1 : n2210_o;
  assign n2212_o = enable_2[77];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2213_o = n1879_o ? 1'b1 : n2212_o;
  assign n2214_o = enable_2[78];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2215_o = n1880_o ? 1'b1 : n2214_o;
  assign n2216_o = enable_2[79];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2217_o = n1881_o ? 1'b1 : n2216_o;
  assign n2218_o = enable_2[80];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2219_o = n1882_o ? 1'b1 : n2218_o;
  assign n2220_o = enable_2[81];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2221_o = n1883_o ? 1'b1 : n2220_o;
  assign n2222_o = enable_2[82];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2223_o = n1884_o ? 1'b1 : n2222_o;
  assign n2224_o = enable_2[83];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2225_o = n1885_o ? 1'b1 : n2224_o;
  assign n2226_o = enable_2[84];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2227_o = n1886_o ? 1'b1 : n2226_o;
  assign n2228_o = enable_2[85];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2229_o = n1887_o ? 1'b1 : n2228_o;
  assign n2230_o = enable_2[86];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2231_o = n1888_o ? 1'b1 : n2230_o;
  assign n2232_o = enable_2[87];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2233_o = n1889_o ? 1'b1 : n2232_o;
  assign n2234_o = enable_2[88];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2235_o = n1890_o ? 1'b1 : n2234_o;
  assign n2236_o = enable_2[89];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2237_o = n1891_o ? 1'b1 : n2236_o;
  assign n2238_o = enable_2[90];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2239_o = n1892_o ? 1'b1 : n2238_o;
  assign n2240_o = enable_2[91];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2241_o = n1893_o ? 1'b1 : n2240_o;
  assign n2242_o = enable_2[92];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2243_o = n1894_o ? 1'b1 : n2242_o;
  assign n2244_o = enable_2[93];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2245_o = n1895_o ? 1'b1 : n2244_o;
  assign n2246_o = enable_2[94];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2247_o = n1896_o ? 1'b1 : n2246_o;
  assign n2248_o = enable_2[95];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2249_o = n1897_o ? 1'b1 : n2248_o;
  assign n2250_o = enable_2[96];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2251_o = n1898_o ? 1'b1 : n2250_o;
  assign n2252_o = enable_2[97];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2253_o = n1899_o ? 1'b1 : n2252_o;
  assign n2254_o = enable_2[98];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2255_o = n1900_o ? 1'b1 : n2254_o;
  assign n2256_o = enable_2[99];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2257_o = n1901_o ? 1'b1 : n2256_o;
  assign n2258_o = enable_2[100];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2259_o = n1902_o ? 1'b1 : n2258_o;
  assign n2260_o = enable_2[101];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2261_o = n1903_o ? 1'b1 : n2260_o;
  assign n2262_o = enable_2[102];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2263_o = n1904_o ? 1'b1 : n2262_o;
  assign n2264_o = enable_2[103];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2265_o = n1905_o ? 1'b1 : n2264_o;
  assign n2266_o = enable_2[104];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2267_o = n1906_o ? 1'b1 : n2266_o;
  assign n2268_o = enable_2[105];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2269_o = n1907_o ? 1'b1 : n2268_o;
  assign n2270_o = enable_2[106];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2271_o = n1908_o ? 1'b1 : n2270_o;
  assign n2272_o = enable_2[107];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2273_o = n1909_o ? 1'b1 : n2272_o;
  assign n2274_o = enable_2[108];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2275_o = n1910_o ? 1'b1 : n2274_o;
  assign n2276_o = enable_2[109];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2277_o = n1911_o ? 1'b1 : n2276_o;
  assign n2278_o = enable_2[110];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2279_o = n1912_o ? 1'b1 : n2278_o;
  assign n2280_o = enable_2[111];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2281_o = n1913_o ? 1'b1 : n2280_o;
  assign n2282_o = enable_2[112];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2283_o = n1914_o ? 1'b1 : n2282_o;
  assign n2284_o = enable_2[113];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2285_o = n1915_o ? 1'b1 : n2284_o;
  assign n2286_o = enable_2[114];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2287_o = n1916_o ? 1'b1 : n2286_o;
  assign n2288_o = enable_2[115];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2289_o = n1917_o ? 1'b1 : n2288_o;
  assign n2290_o = enable_2[116];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2291_o = n1918_o ? 1'b1 : n2290_o;
  assign n2292_o = enable_2[117];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2293_o = n1919_o ? 1'b1 : n2292_o;
  assign n2294_o = enable_2[118];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2295_o = n1920_o ? 1'b1 : n2294_o;
  assign n2296_o = enable_2[119];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2297_o = n1921_o ? 1'b1 : n2296_o;
  assign n2298_o = enable_2[120];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2299_o = n1922_o ? 1'b1 : n2298_o;
  assign n2300_o = enable_2[121];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2301_o = n1923_o ? 1'b1 : n2300_o;
  assign n2302_o = enable_2[122];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2303_o = n1924_o ? 1'b1 : n2302_o;
  assign n2304_o = enable_2[123];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2305_o = n1925_o ? 1'b1 : n2304_o;
  assign n2306_o = enable_2[124];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2307_o = n1926_o ? 1'b1 : n2306_o;
  assign n2308_o = enable_2[125];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2309_o = n1927_o ? 1'b1 : n2308_o;
  assign n2310_o = enable_2[126];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2311_o = n1928_o ? 1'b1 : n2310_o;
  assign n2312_o = enable_2[127];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2313_o = n1929_o ? 1'b1 : n2312_o;
  assign n2314_o = enable_2[128];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2315_o = n1930_o ? 1'b1 : n2314_o;
  assign n2316_o = enable_2[129];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2317_o = n1931_o ? 1'b1 : n2316_o;
  assign n2318_o = enable_2[130];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2319_o = n1932_o ? 1'b1 : n2318_o;
  assign n2320_o = enable_2[131];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2321_o = n1933_o ? 1'b1 : n2320_o;
  assign n2322_o = enable_2[132];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2323_o = n1934_o ? 1'b1 : n2322_o;
  assign n2324_o = enable_2[133];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2325_o = n1935_o ? 1'b1 : n2324_o;
  assign n2326_o = enable_2[134];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2327_o = n1936_o ? 1'b1 : n2326_o;
  assign n2328_o = enable_2[135];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2329_o = n1937_o ? 1'b1 : n2328_o;
  assign n2330_o = enable_2[136];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2331_o = n1938_o ? 1'b1 : n2330_o;
  assign n2332_o = enable_2[137];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2333_o = n1939_o ? 1'b1 : n2332_o;
  assign n2334_o = enable_2[138];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2335_o = n1940_o ? 1'b1 : n2334_o;
  assign n2336_o = enable_2[139];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2337_o = n1941_o ? 1'b1 : n2336_o;
  assign n2338_o = enable_2[140];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2339_o = n1942_o ? 1'b1 : n2338_o;
  assign n2340_o = enable_2[141];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2341_o = n1943_o ? 1'b1 : n2340_o;
  assign n2342_o = enable_2[142];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2343_o = n1944_o ? 1'b1 : n2342_o;
  assign n2344_o = enable_2[143];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2345_o = n1945_o ? 1'b1 : n2344_o;
  assign n2346_o = enable_2[144];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2347_o = n1946_o ? 1'b1 : n2346_o;
  assign n2348_o = enable_2[145];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2349_o = n1947_o ? 1'b1 : n2348_o;
  assign n2350_o = enable_2[146];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2351_o = n1948_o ? 1'b1 : n2350_o;
  assign n2352_o = enable_2[147];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2353_o = n1949_o ? 1'b1 : n2352_o;
  assign n2354_o = enable_2[148];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2355_o = n1950_o ? 1'b1 : n2354_o;
  assign n2356_o = enable_2[149];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2357_o = n1951_o ? 1'b1 : n2356_o;
  assign n2358_o = enable_2[150];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2359_o = n1952_o ? 1'b1 : n2358_o;
  assign n2360_o = enable_2[151];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2361_o = n1953_o ? 1'b1 : n2360_o;
  assign n2362_o = enable_2[152];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2363_o = n1954_o ? 1'b1 : n2362_o;
  assign n2364_o = enable_2[153];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2365_o = n1955_o ? 1'b1 : n2364_o;
  assign n2366_o = enable_2[154];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2367_o = n1956_o ? 1'b1 : n2366_o;
  assign n2368_o = enable_2[155];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2369_o = n1957_o ? 1'b1 : n2368_o;
  assign n2370_o = enable_2[156];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2371_o = n1958_o ? 1'b1 : n2370_o;
  assign n2372_o = enable_2[157];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2373_o = n1959_o ? 1'b1 : n2372_o;
  assign n2374_o = enable_2[158];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2375_o = n1960_o ? 1'b1 : n2374_o;
  assign n2376_o = enable_2[159];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2377_o = n1961_o ? 1'b1 : n2376_o;
  assign n2378_o = enable_2[160];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2379_o = n1962_o ? 1'b1 : n2378_o;
  assign n2380_o = enable_2[161];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2381_o = n1963_o ? 1'b1 : n2380_o;
  assign n2382_o = enable_2[162];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2383_o = n1964_o ? 1'b1 : n2382_o;
  assign n2384_o = enable_2[163];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2385_o = n1965_o ? 1'b1 : n2384_o;
  assign n2386_o = enable_2[164];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2387_o = n1966_o ? 1'b1 : n2386_o;
  assign n2388_o = enable_2[165];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2389_o = n1967_o ? 1'b1 : n2388_o;
  assign n2390_o = enable_2[166];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2391_o = n1968_o ? 1'b1 : n2390_o;
  assign n2392_o = enable_2[167];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2393_o = n1969_o ? 1'b1 : n2392_o;
  assign n2394_o = enable_2[168];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2395_o = n1970_o ? 1'b1 : n2394_o;
  assign n2396_o = enable_2[169];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2397_o = n1971_o ? 1'b1 : n2396_o;
  assign n2398_o = enable_2[170];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2399_o = n1972_o ? 1'b1 : n2398_o;
  assign n2400_o = enable_2[171];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2401_o = n1973_o ? 1'b1 : n2400_o;
  assign n2402_o = enable_2[172];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2403_o = n1974_o ? 1'b1 : n2402_o;
  assign n2404_o = enable_2[173];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2405_o = n1975_o ? 1'b1 : n2404_o;
  assign n2406_o = enable_2[174];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2407_o = n1976_o ? 1'b1 : n2406_o;
  assign n2408_o = enable_2[175];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2409_o = n1977_o ? 1'b1 : n2408_o;
  assign n2410_o = enable_2[176];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2411_o = n1978_o ? 1'b1 : n2410_o;
  assign n2412_o = enable_2[177];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2413_o = n1979_o ? 1'b1 : n2412_o;
  assign n2414_o = enable_2[178];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2415_o = n1980_o ? 1'b1 : n2414_o;
  assign n2416_o = enable_2[179];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2417_o = n1981_o ? 1'b1 : n2416_o;
  assign n2418_o = enable_2[180];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2419_o = n1982_o ? 1'b1 : n2418_o;
  assign n2420_o = enable_2[181];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2421_o = n1983_o ? 1'b1 : n2420_o;
  assign n2422_o = enable_2[182];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2423_o = n1984_o ? 1'b1 : n2422_o;
  assign n2424_o = enable_2[183];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2425_o = n1985_o ? 1'b1 : n2424_o;
  assign n2426_o = enable_2[184];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2427_o = n1986_o ? 1'b1 : n2426_o;
  assign n2428_o = enable_2[185];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2429_o = n1987_o ? 1'b1 : n2428_o;
  assign n2430_o = enable_2[186];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2431_o = n1988_o ? 1'b1 : n2430_o;
  assign n2432_o = enable_2[187];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2433_o = n1989_o ? 1'b1 : n2432_o;
  assign n2434_o = enable_2[188];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2435_o = n1990_o ? 1'b1 : n2434_o;
  assign n2436_o = enable_2[189];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2437_o = n1991_o ? 1'b1 : n2436_o;
  assign n2438_o = enable_2[190];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2439_o = n1992_o ? 1'b1 : n2438_o;
  assign n2440_o = enable_2[191];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2441_o = n1993_o ? 1'b1 : n2440_o;
  assign n2442_o = enable_2[192];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2443_o = n1994_o ? 1'b1 : n2442_o;
  assign n2444_o = enable_2[193];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2445_o = n1995_o ? 1'b1 : n2444_o;
  assign n2446_o = enable_2[194];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2447_o = n1996_o ? 1'b1 : n2446_o;
  assign n2448_o = enable_2[195];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2449_o = n1997_o ? 1'b1 : n2448_o;
  assign n2450_o = enable_2[196];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2451_o = n1998_o ? 1'b1 : n2450_o;
  assign n2452_o = enable_2[197];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2453_o = n1999_o ? 1'b1 : n2452_o;
  assign n2454_o = enable_2[198];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2455_o = n2000_o ? 1'b1 : n2454_o;
  assign n2456_o = enable_2[199];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2457_o = n2001_o ? 1'b1 : n2456_o;
  assign n2458_o = enable_2[200];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2459_o = n2002_o ? 1'b1 : n2458_o;
  assign n2460_o = enable_2[201];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2461_o = n2003_o ? 1'b1 : n2460_o;
  assign n2462_o = enable_2[202];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2463_o = n2004_o ? 1'b1 : n2462_o;
  assign n2464_o = enable_2[203];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2465_o = n2005_o ? 1'b1 : n2464_o;
  assign n2466_o = enable_2[204];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2467_o = n2006_o ? 1'b1 : n2466_o;
  assign n2468_o = enable_2[205];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2469_o = n2007_o ? 1'b1 : n2468_o;
  assign n2470_o = enable_2[206];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2471_o = n2008_o ? 1'b1 : n2470_o;
  assign n2472_o = enable_2[207];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2473_o = n2009_o ? 1'b1 : n2472_o;
  assign n2474_o = enable_2[208];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2475_o = n2010_o ? 1'b1 : n2474_o;
  assign n2476_o = enable_2[209];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2477_o = n2011_o ? 1'b1 : n2476_o;
  assign n2478_o = enable_2[210];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2479_o = n2012_o ? 1'b1 : n2478_o;
  assign n2480_o = enable_2[211];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2481_o = n2013_o ? 1'b1 : n2480_o;
  assign n2482_o = enable_2[212];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2483_o = n2014_o ? 1'b1 : n2482_o;
  assign n2484_o = enable_2[213];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2485_o = n2015_o ? 1'b1 : n2484_o;
  assign n2486_o = enable_2[214];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2487_o = n2016_o ? 1'b1 : n2486_o;
  assign n2488_o = enable_2[215];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2489_o = n2017_o ? 1'b1 : n2488_o;
  assign n2490_o = enable_2[216];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2491_o = n2018_o ? 1'b1 : n2490_o;
  assign n2492_o = enable_2[217];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2493_o = n2019_o ? 1'b1 : n2492_o;
  assign n2494_o = enable_2[218];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2495_o = n2020_o ? 1'b1 : n2494_o;
  assign n2496_o = enable_2[219];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2497_o = n2021_o ? 1'b1 : n2496_o;
  assign n2498_o = enable_2[220];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2499_o = n2022_o ? 1'b1 : n2498_o;
  assign n2500_o = enable_2[221];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2501_o = n2023_o ? 1'b1 : n2500_o;
  assign n2502_o = enable_2[222];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2503_o = n2024_o ? 1'b1 : n2502_o;
  assign n2504_o = enable_2[223];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2505_o = n2025_o ? 1'b1 : n2504_o;
  assign n2506_o = enable_2[224];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2507_o = n2026_o ? 1'b1 : n2506_o;
  assign n2508_o = enable_2[225];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2509_o = n2027_o ? 1'b1 : n2508_o;
  assign n2510_o = enable_2[226];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2511_o = n2028_o ? 1'b1 : n2510_o;
  assign n2512_o = enable_2[227];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2513_o = n2029_o ? 1'b1 : n2512_o;
  assign n2514_o = enable_2[228];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2515_o = n2030_o ? 1'b1 : n2514_o;
  assign n2516_o = enable_2[229];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2517_o = n2031_o ? 1'b1 : n2516_o;
  assign n2518_o = enable_2[230];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2519_o = n2032_o ? 1'b1 : n2518_o;
  assign n2520_o = enable_2[231];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2521_o = n2033_o ? 1'b1 : n2520_o;
  assign n2522_o = enable_2[232];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2523_o = n2034_o ? 1'b1 : n2522_o;
  assign n2524_o = enable_2[233];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2525_o = n2035_o ? 1'b1 : n2524_o;
  assign n2526_o = enable_2[234];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2527_o = n2036_o ? 1'b1 : n2526_o;
  assign n2528_o = enable_2[235];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2529_o = n2037_o ? 1'b1 : n2528_o;
  assign n2530_o = enable_2[236];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2531_o = n2038_o ? 1'b1 : n2530_o;
  assign n2532_o = enable_2[237];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2533_o = n2039_o ? 1'b1 : n2532_o;
  assign n2534_o = enable_2[238];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2535_o = n2040_o ? 1'b1 : n2534_o;
  assign n2536_o = enable_2[239];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2537_o = n2041_o ? 1'b1 : n2536_o;
  assign n2538_o = enable_2[240];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2539_o = n2042_o ? 1'b1 : n2538_o;
  assign n2540_o = enable_2[241];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2541_o = n2043_o ? 1'b1 : n2540_o;
  assign n2542_o = enable_2[242];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2543_o = n2044_o ? 1'b1 : n2542_o;
  assign n2544_o = enable_2[243];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2545_o = n2045_o ? 1'b1 : n2544_o;
  assign n2546_o = enable_2[244];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2547_o = n2046_o ? 1'b1 : n2546_o;
  assign n2548_o = enable_2[245];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2549_o = n2047_o ? 1'b1 : n2548_o;
  assign n2550_o = enable_2[246];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2551_o = n2048_o ? 1'b1 : n2550_o;
  assign n2552_o = enable_2[247];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2553_o = n2049_o ? 1'b1 : n2552_o;
  assign n2554_o = enable_2[248];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2555_o = n2050_o ? 1'b1 : n2554_o;
  assign n2556_o = enable_2[249];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2557_o = n2051_o ? 1'b1 : n2556_o;
  assign n2558_o = enable_2[250];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2559_o = n2052_o ? 1'b1 : n2558_o;
  assign n2560_o = enable_2[251];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2561_o = n2053_o ? 1'b1 : n2560_o;
  assign n2562_o = enable_2[252];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2563_o = n2054_o ? 1'b1 : n2562_o;
  assign n2564_o = enable_2[253];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2565_o = n2055_o ? 1'b1 : n2564_o;
  assign n2566_o = enable_2[254];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2567_o = n2056_o ? 1'b1 : n2566_o;
  assign n2568_o = enable_2[255];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:435:21  */
  assign n2569_o = n2057_o ? 1'b1 : n2568_o;
  assign n2570_o = {n2569_o, n2567_o, n2565_o, n2563_o, n2561_o, n2559_o, n2557_o, n2555_o, n2553_o, n2551_o, n2549_o, n2547_o, n2545_o, n2543_o, n2541_o, n2539_o, n2537_o, n2535_o, n2533_o, n2531_o, n2529_o, n2527_o, n2525_o, n2523_o, n2521_o, n2519_o, n2517_o, n2515_o, n2513_o, n2511_o, n2509_o, n2507_o, n2505_o, n2503_o, n2501_o, n2499_o, n2497_o, n2495_o, n2493_o, n2491_o, n2489_o, n2487_o, n2485_o, n2483_o, n2481_o, n2479_o, n2477_o, n2475_o, n2473_o, n2471_o, n2469_o, n2467_o, n2465_o, n2463_o, n2461_o, n2459_o, n2457_o, n2455_o, n2453_o, n2451_o, n2449_o, n2447_o, n2445_o, n2443_o, n2441_o, n2439_o, n2437_o, n2435_o, n2433_o, n2431_o, n2429_o, n2427_o, n2425_o, n2423_o, n2421_o, n2419_o, n2417_o, n2415_o, n2413_o, n2411_o, n2409_o, n2407_o, n2405_o, n2403_o, n2401_o, n2399_o, n2397_o, n2395_o, n2393_o, n2391_o, n2389_o, n2387_o, n2385_o, n2383_o, n2381_o, n2379_o, n2377_o, n2375_o, n2373_o, n2371_o, n2369_o, n2367_o, n2365_o, n2363_o, n2361_o, n2359_o, n2357_o, n2355_o, n2353_o, n2351_o, n2349_o, n2347_o, n2345_o, n2343_o, n2341_o, n2339_o, n2337_o, n2335_o, n2333_o, n2331_o, n2329_o, n2327_o, n2325_o, n2323_o, n2321_o, n2319_o, n2317_o, n2315_o, n2313_o, n2311_o, n2309_o, n2307_o, n2305_o, n2303_o, n2301_o, n2299_o, n2297_o, n2295_o, n2293_o, n2291_o, n2289_o, n2287_o, n2285_o, n2283_o, n2281_o, n2279_o, n2277_o, n2275_o, n2273_o, n2271_o, n2269_o, n2267_o, n2265_o, n2263_o, n2261_o, n2259_o, n2257_o, n2255_o, n2253_o, n2251_o, n2249_o, n2247_o, n2245_o, n2243_o, n2241_o, n2239_o, n2237_o, n2235_o, n2233_o, n2231_o, n2229_o, n2227_o, n2225_o, n2223_o, n2221_o, n2219_o, n2217_o, n2215_o, n2213_o, n2211_o, n2209_o, n2207_o, n2205_o, n2203_o, n2201_o, n2199_o, n2197_o, n2195_o, n2193_o, n2191_o, n2189_o, n2187_o, n2185_o, n2183_o, n2181_o, n2179_o, n2177_o, n2175_o, n2173_o, n2171_o, n2169_o, n2167_o, n2165_o, n2163_o, n2161_o, n2159_o, n2157_o, n2155_o, n2153_o, n2151_o, n2149_o, n2147_o, n2145_o, n2143_o, n2141_o, n2139_o, n2137_o, n2135_o, n2133_o, n2131_o, n2129_o, n2127_o, n2125_o, n2123_o, n2121_o, n2119_o, n2117_o, n2115_o, n2113_o, n2111_o, n2109_o, n2107_o, n2105_o, n2103_o, n2101_o, n2099_o, n2097_o, n2095_o, n2093_o, n2091_o, n2089_o, n2087_o, n2085_o, n2083_o, n2081_o, n2079_o, n2077_o, n2075_o, n2073_o, n2071_o, n2069_o, n2067_o, n2065_o, n2063_o, n2061_o, n2059_o};
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2571_o = n262_o[7];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2572_o = ~n2571_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2573_o = n262_o[6];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2574_o = ~n2573_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2575_o = n2572_o & n2574_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2576_o = n2572_o & n2573_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2577_o = n2571_o & n2574_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2578_o = n2571_o & n2573_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2579_o = n262_o[5];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2580_o = ~n2579_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2581_o = n2575_o & n2580_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2582_o = n2575_o & n2579_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2583_o = n2576_o & n2580_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2584_o = n2576_o & n2579_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2585_o = n2577_o & n2580_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2586_o = n2577_o & n2579_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2587_o = n2578_o & n2580_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2588_o = n2578_o & n2579_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2589_o = n262_o[4];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2590_o = ~n2589_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2591_o = n2581_o & n2590_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2592_o = n2581_o & n2589_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2593_o = n2582_o & n2590_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2594_o = n2582_o & n2589_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2595_o = n2583_o & n2590_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2596_o = n2583_o & n2589_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2597_o = n2584_o & n2590_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2598_o = n2584_o & n2589_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2599_o = n2585_o & n2590_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2600_o = n2585_o & n2589_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2601_o = n2586_o & n2590_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2602_o = n2586_o & n2589_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2603_o = n2587_o & n2590_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2604_o = n2587_o & n2589_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2605_o = n2588_o & n2590_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2606_o = n2588_o & n2589_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2607_o = n262_o[3];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2608_o = ~n2607_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2609_o = n2591_o & n2608_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2610_o = n2591_o & n2607_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2611_o = n2592_o & n2608_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2612_o = n2592_o & n2607_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2613_o = n2593_o & n2608_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2614_o = n2593_o & n2607_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2615_o = n2594_o & n2608_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2616_o = n2594_o & n2607_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2617_o = n2595_o & n2608_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2618_o = n2595_o & n2607_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2619_o = n2596_o & n2608_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2620_o = n2596_o & n2607_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2621_o = n2597_o & n2608_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2622_o = n2597_o & n2607_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2623_o = n2598_o & n2608_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2624_o = n2598_o & n2607_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2625_o = n2599_o & n2608_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2626_o = n2599_o & n2607_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2627_o = n2600_o & n2608_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2628_o = n2600_o & n2607_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2629_o = n2601_o & n2608_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2630_o = n2601_o & n2607_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2631_o = n2602_o & n2608_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2632_o = n2602_o & n2607_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2633_o = n2603_o & n2608_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2634_o = n2603_o & n2607_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2635_o = n2604_o & n2608_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2636_o = n2604_o & n2607_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2637_o = n2605_o & n2608_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2638_o = n2605_o & n2607_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2639_o = n2606_o & n2608_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2640_o = n2606_o & n2607_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2641_o = n262_o[2];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2642_o = ~n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2643_o = n2609_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2644_o = n2609_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2645_o = n2610_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2646_o = n2610_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2647_o = n2611_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2648_o = n2611_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2649_o = n2612_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2650_o = n2612_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2651_o = n2613_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2652_o = n2613_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2653_o = n2614_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2654_o = n2614_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2655_o = n2615_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2656_o = n2615_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2657_o = n2616_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2658_o = n2616_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2659_o = n2617_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2660_o = n2617_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2661_o = n2618_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2662_o = n2618_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2663_o = n2619_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2664_o = n2619_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2665_o = n2620_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2666_o = n2620_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2667_o = n2621_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2668_o = n2621_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2669_o = n2622_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2670_o = n2622_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2671_o = n2623_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2672_o = n2623_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2673_o = n2624_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2674_o = n2624_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2675_o = n2625_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2676_o = n2625_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2677_o = n2626_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2678_o = n2626_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2679_o = n2627_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2680_o = n2627_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2681_o = n2628_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2682_o = n2628_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2683_o = n2629_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2684_o = n2629_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2685_o = n2630_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2686_o = n2630_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2687_o = n2631_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2688_o = n2631_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2689_o = n2632_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2690_o = n2632_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2691_o = n2633_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2692_o = n2633_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2693_o = n2634_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2694_o = n2634_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2695_o = n2635_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2696_o = n2635_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2697_o = n2636_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2698_o = n2636_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2699_o = n2637_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2700_o = n2637_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2701_o = n2638_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2702_o = n2638_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2703_o = n2639_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2704_o = n2639_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2705_o = n2640_o & n2642_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2706_o = n2640_o & n2641_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2707_o = n262_o[1];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2708_o = ~n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2709_o = n2643_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2710_o = n2643_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2711_o = n2644_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2712_o = n2644_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2713_o = n2645_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2714_o = n2645_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2715_o = n2646_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2716_o = n2646_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2717_o = n2647_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2718_o = n2647_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2719_o = n2648_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2720_o = n2648_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2721_o = n2649_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2722_o = n2649_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2723_o = n2650_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2724_o = n2650_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2725_o = n2651_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2726_o = n2651_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2727_o = n2652_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2728_o = n2652_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2729_o = n2653_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2730_o = n2653_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2731_o = n2654_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2732_o = n2654_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2733_o = n2655_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2734_o = n2655_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2735_o = n2656_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2736_o = n2656_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2737_o = n2657_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2738_o = n2657_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2739_o = n2658_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2740_o = n2658_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2741_o = n2659_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2742_o = n2659_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2743_o = n2660_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2744_o = n2660_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2745_o = n2661_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2746_o = n2661_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2747_o = n2662_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2748_o = n2662_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2749_o = n2663_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2750_o = n2663_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2751_o = n2664_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2752_o = n2664_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2753_o = n2665_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2754_o = n2665_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2755_o = n2666_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2756_o = n2666_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2757_o = n2667_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2758_o = n2667_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2759_o = n2668_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2760_o = n2668_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2761_o = n2669_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2762_o = n2669_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2763_o = n2670_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2764_o = n2670_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2765_o = n2671_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2766_o = n2671_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2767_o = n2672_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2768_o = n2672_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2769_o = n2673_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2770_o = n2673_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2771_o = n2674_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2772_o = n2674_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2773_o = n2675_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2774_o = n2675_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2775_o = n2676_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2776_o = n2676_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2777_o = n2677_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2778_o = n2677_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2779_o = n2678_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2780_o = n2678_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2781_o = n2679_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2782_o = n2679_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2783_o = n2680_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2784_o = n2680_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2785_o = n2681_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2786_o = n2681_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2787_o = n2682_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2788_o = n2682_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2789_o = n2683_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2790_o = n2683_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2791_o = n2684_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2792_o = n2684_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2793_o = n2685_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2794_o = n2685_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2795_o = n2686_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2796_o = n2686_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2797_o = n2687_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2798_o = n2687_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2799_o = n2688_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2800_o = n2688_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2801_o = n2689_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2802_o = n2689_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2803_o = n2690_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2804_o = n2690_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2805_o = n2691_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2806_o = n2691_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2807_o = n2692_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2808_o = n2692_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2809_o = n2693_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2810_o = n2693_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2811_o = n2694_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2812_o = n2694_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2813_o = n2695_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2814_o = n2695_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2815_o = n2696_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2816_o = n2696_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2817_o = n2697_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2818_o = n2697_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2819_o = n2698_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2820_o = n2698_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2821_o = n2699_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2822_o = n2699_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2823_o = n2700_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2824_o = n2700_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2825_o = n2701_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2826_o = n2701_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2827_o = n2702_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2828_o = n2702_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2829_o = n2703_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2830_o = n2703_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2831_o = n2704_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2832_o = n2704_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2833_o = n2705_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2834_o = n2705_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2835_o = n2706_o & n2708_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2836_o = n2706_o & n2707_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2837_o = n262_o[0];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2838_o = ~n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2839_o = n2709_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2840_o = n2709_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2841_o = n2710_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2842_o = n2710_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2843_o = n2711_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2844_o = n2711_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2845_o = n2712_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2846_o = n2712_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2847_o = n2713_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2848_o = n2713_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2849_o = n2714_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2850_o = n2714_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2851_o = n2715_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2852_o = n2715_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2853_o = n2716_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2854_o = n2716_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2855_o = n2717_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2856_o = n2717_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2857_o = n2718_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2858_o = n2718_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2859_o = n2719_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2860_o = n2719_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2861_o = n2720_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2862_o = n2720_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2863_o = n2721_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2864_o = n2721_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2865_o = n2722_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2866_o = n2722_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2867_o = n2723_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2868_o = n2723_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2869_o = n2724_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2870_o = n2724_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2871_o = n2725_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2872_o = n2725_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2873_o = n2726_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2874_o = n2726_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2875_o = n2727_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2876_o = n2727_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2877_o = n2728_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2878_o = n2728_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2879_o = n2729_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2880_o = n2729_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2881_o = n2730_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2882_o = n2730_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2883_o = n2731_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2884_o = n2731_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2885_o = n2732_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2886_o = n2732_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2887_o = n2733_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2888_o = n2733_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2889_o = n2734_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2890_o = n2734_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2891_o = n2735_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2892_o = n2735_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2893_o = n2736_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2894_o = n2736_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2895_o = n2737_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2896_o = n2737_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2897_o = n2738_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2898_o = n2738_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2899_o = n2739_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2900_o = n2739_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2901_o = n2740_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2902_o = n2740_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2903_o = n2741_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2904_o = n2741_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2905_o = n2742_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2906_o = n2742_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2907_o = n2743_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2908_o = n2743_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2909_o = n2744_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2910_o = n2744_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2911_o = n2745_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2912_o = n2745_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2913_o = n2746_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2914_o = n2746_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2915_o = n2747_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2916_o = n2747_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2917_o = n2748_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2918_o = n2748_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2919_o = n2749_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2920_o = n2749_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2921_o = n2750_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2922_o = n2750_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2923_o = n2751_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2924_o = n2751_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2925_o = n2752_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2926_o = n2752_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2927_o = n2753_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2928_o = n2753_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2929_o = n2754_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2930_o = n2754_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2931_o = n2755_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2932_o = n2755_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2933_o = n2756_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2934_o = n2756_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2935_o = n2757_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2936_o = n2757_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2937_o = n2758_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2938_o = n2758_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2939_o = n2759_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2940_o = n2759_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2941_o = n2760_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2942_o = n2760_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2943_o = n2761_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2944_o = n2761_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2945_o = n2762_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2946_o = n2762_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2947_o = n2763_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2948_o = n2763_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2949_o = n2764_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2950_o = n2764_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2951_o = n2765_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2952_o = n2765_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2953_o = n2766_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2954_o = n2766_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2955_o = n2767_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2956_o = n2767_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2957_o = n2768_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2958_o = n2768_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2959_o = n2769_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2960_o = n2769_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2961_o = n2770_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2962_o = n2770_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2963_o = n2771_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2964_o = n2771_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2965_o = n2772_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2966_o = n2772_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2967_o = n2773_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2968_o = n2773_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2969_o = n2774_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2970_o = n2774_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2971_o = n2775_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2972_o = n2775_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2973_o = n2776_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2974_o = n2776_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2975_o = n2777_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2976_o = n2777_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2977_o = n2778_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2978_o = n2778_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2979_o = n2779_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2980_o = n2779_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2981_o = n2780_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2982_o = n2780_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2983_o = n2781_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2984_o = n2781_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2985_o = n2782_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2986_o = n2782_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2987_o = n2783_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2988_o = n2783_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2989_o = n2784_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2990_o = n2784_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2991_o = n2785_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2992_o = n2785_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2993_o = n2786_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2994_o = n2786_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2995_o = n2787_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2996_o = n2787_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2997_o = n2788_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2998_o = n2788_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n2999_o = n2789_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3000_o = n2789_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3001_o = n2790_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3002_o = n2790_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3003_o = n2791_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3004_o = n2791_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3005_o = n2792_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3006_o = n2792_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3007_o = n2793_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3008_o = n2793_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3009_o = n2794_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3010_o = n2794_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3011_o = n2795_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3012_o = n2795_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3013_o = n2796_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3014_o = n2796_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3015_o = n2797_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3016_o = n2797_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3017_o = n2798_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3018_o = n2798_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3019_o = n2799_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3020_o = n2799_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3021_o = n2800_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3022_o = n2800_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3023_o = n2801_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3024_o = n2801_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3025_o = n2802_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3026_o = n2802_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3027_o = n2803_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3028_o = n2803_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3029_o = n2804_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3030_o = n2804_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3031_o = n2805_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3032_o = n2805_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3033_o = n2806_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3034_o = n2806_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3035_o = n2807_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3036_o = n2807_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3037_o = n2808_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3038_o = n2808_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3039_o = n2809_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3040_o = n2809_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3041_o = n2810_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3042_o = n2810_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3043_o = n2811_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3044_o = n2811_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3045_o = n2812_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3046_o = n2812_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3047_o = n2813_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3048_o = n2813_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3049_o = n2814_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3050_o = n2814_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3051_o = n2815_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3052_o = n2815_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3053_o = n2816_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3054_o = n2816_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3055_o = n2817_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3056_o = n2817_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3057_o = n2818_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3058_o = n2818_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3059_o = n2819_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3060_o = n2819_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3061_o = n2820_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3062_o = n2820_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3063_o = n2821_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3064_o = n2821_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3065_o = n2822_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3066_o = n2822_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3067_o = n2823_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3068_o = n2823_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3069_o = n2824_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3070_o = n2824_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3071_o = n2825_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3072_o = n2825_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3073_o = n2826_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3074_o = n2826_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3075_o = n2827_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3076_o = n2827_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3077_o = n2828_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3078_o = n2828_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3079_o = n2829_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3080_o = n2829_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3081_o = n2830_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3082_o = n2830_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3083_o = n2831_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3084_o = n2831_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3085_o = n2832_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3086_o = n2832_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3087_o = n2833_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3088_o = n2833_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3089_o = n2834_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3090_o = n2834_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3091_o = n2835_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3092_o = n2835_o & n2837_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3093_o = n2836_o & n2838_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3094_o = n2836_o & n2837_o;
  assign n3095_o = enable_1[0];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3096_o = n2839_o ? 1'b1 : n3095_o;
  assign n3097_o = enable_1[1];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3098_o = n2840_o ? 1'b1 : n3097_o;
  assign n3099_o = enable_1[2];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3100_o = n2841_o ? 1'b1 : n3099_o;
  assign n3101_o = enable_1[3];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3102_o = n2842_o ? 1'b1 : n3101_o;
  assign n3103_o = enable_1[4];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3104_o = n2843_o ? 1'b1 : n3103_o;
  assign n3105_o = enable_1[5];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3106_o = n2844_o ? 1'b1 : n3105_o;
  assign n3107_o = enable_1[6];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3108_o = n2845_o ? 1'b1 : n3107_o;
  assign n3109_o = enable_1[7];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3110_o = n2846_o ? 1'b1 : n3109_o;
  assign n3111_o = enable_1[8];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3112_o = n2847_o ? 1'b1 : n3111_o;
  assign n3113_o = enable_1[9];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3114_o = n2848_o ? 1'b1 : n3113_o;
  assign n3115_o = enable_1[10];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3116_o = n2849_o ? 1'b1 : n3115_o;
  assign n3117_o = enable_1[11];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3118_o = n2850_o ? 1'b1 : n3117_o;
  assign n3119_o = enable_1[12];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3120_o = n2851_o ? 1'b1 : n3119_o;
  assign n3121_o = enable_1[13];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3122_o = n2852_o ? 1'b1 : n3121_o;
  assign n3123_o = enable_1[14];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3124_o = n2853_o ? 1'b1 : n3123_o;
  assign n3125_o = enable_1[15];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3126_o = n2854_o ? 1'b1 : n3125_o;
  assign n3127_o = enable_1[16];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3128_o = n2855_o ? 1'b1 : n3127_o;
  assign n3129_o = enable_1[17];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3130_o = n2856_o ? 1'b1 : n3129_o;
  assign n3131_o = enable_1[18];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3132_o = n2857_o ? 1'b1 : n3131_o;
  assign n3133_o = enable_1[19];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3134_o = n2858_o ? 1'b1 : n3133_o;
  assign n3135_o = enable_1[20];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3136_o = n2859_o ? 1'b1 : n3135_o;
  assign n3137_o = enable_1[21];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3138_o = n2860_o ? 1'b1 : n3137_o;
  assign n3139_o = enable_1[22];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3140_o = n2861_o ? 1'b1 : n3139_o;
  assign n3141_o = enable_1[23];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3142_o = n2862_o ? 1'b1 : n3141_o;
  assign n3143_o = enable_1[24];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3144_o = n2863_o ? 1'b1 : n3143_o;
  assign n3145_o = enable_1[25];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3146_o = n2864_o ? 1'b1 : n3145_o;
  assign n3147_o = enable_1[26];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3148_o = n2865_o ? 1'b1 : n3147_o;
  assign n3149_o = enable_1[27];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3150_o = n2866_o ? 1'b1 : n3149_o;
  assign n3151_o = enable_1[28];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3152_o = n2867_o ? 1'b1 : n3151_o;
  assign n3153_o = enable_1[29];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3154_o = n2868_o ? 1'b1 : n3153_o;
  assign n3155_o = enable_1[30];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3156_o = n2869_o ? 1'b1 : n3155_o;
  assign n3157_o = enable_1[31];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3158_o = n2870_o ? 1'b1 : n3157_o;
  assign n3159_o = enable_1[32];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3160_o = n2871_o ? 1'b1 : n3159_o;
  assign n3161_o = enable_1[33];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3162_o = n2872_o ? 1'b1 : n3161_o;
  assign n3163_o = enable_1[34];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3164_o = n2873_o ? 1'b1 : n3163_o;
  assign n3165_o = enable_1[35];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3166_o = n2874_o ? 1'b1 : n3165_o;
  assign n3167_o = enable_1[36];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3168_o = n2875_o ? 1'b1 : n3167_o;
  assign n3169_o = enable_1[37];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3170_o = n2876_o ? 1'b1 : n3169_o;
  assign n3171_o = enable_1[38];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3172_o = n2877_o ? 1'b1 : n3171_o;
  assign n3173_o = enable_1[39];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3174_o = n2878_o ? 1'b1 : n3173_o;
  assign n3175_o = enable_1[40];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3176_o = n2879_o ? 1'b1 : n3175_o;
  assign n3177_o = enable_1[41];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3178_o = n2880_o ? 1'b1 : n3177_o;
  assign n3179_o = enable_1[42];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3180_o = n2881_o ? 1'b1 : n3179_o;
  assign n3181_o = enable_1[43];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3182_o = n2882_o ? 1'b1 : n3181_o;
  assign n3183_o = enable_1[44];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3184_o = n2883_o ? 1'b1 : n3183_o;
  assign n3185_o = enable_1[45];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3186_o = n2884_o ? 1'b1 : n3185_o;
  assign n3187_o = enable_1[46];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3188_o = n2885_o ? 1'b1 : n3187_o;
  assign n3189_o = enable_1[47];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3190_o = n2886_o ? 1'b1 : n3189_o;
  assign n3191_o = enable_1[48];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3192_o = n2887_o ? 1'b1 : n3191_o;
  assign n3193_o = enable_1[49];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3194_o = n2888_o ? 1'b1 : n3193_o;
  assign n3195_o = enable_1[50];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3196_o = n2889_o ? 1'b1 : n3195_o;
  assign n3197_o = enable_1[51];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3198_o = n2890_o ? 1'b1 : n3197_o;
  assign n3199_o = enable_1[52];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3200_o = n2891_o ? 1'b1 : n3199_o;
  assign n3201_o = enable_1[53];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3202_o = n2892_o ? 1'b1 : n3201_o;
  assign n3203_o = enable_1[54];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3204_o = n2893_o ? 1'b1 : n3203_o;
  assign n3205_o = enable_1[55];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3206_o = n2894_o ? 1'b1 : n3205_o;
  assign n3207_o = enable_1[56];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3208_o = n2895_o ? 1'b1 : n3207_o;
  assign n3209_o = enable_1[57];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3210_o = n2896_o ? 1'b1 : n3209_o;
  assign n3211_o = enable_1[58];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3212_o = n2897_o ? 1'b1 : n3211_o;
  assign n3213_o = enable_1[59];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3214_o = n2898_o ? 1'b1 : n3213_o;
  assign n3215_o = enable_1[60];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3216_o = n2899_o ? 1'b1 : n3215_o;
  assign n3217_o = enable_1[61];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3218_o = n2900_o ? 1'b1 : n3217_o;
  assign n3219_o = enable_1[62];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3220_o = n2901_o ? 1'b1 : n3219_o;
  assign n3221_o = enable_1[63];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3222_o = n2902_o ? 1'b1 : n3221_o;
  assign n3223_o = enable_1[64];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3224_o = n2903_o ? 1'b1 : n3223_o;
  assign n3225_o = enable_1[65];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3226_o = n2904_o ? 1'b1 : n3225_o;
  assign n3227_o = enable_1[66];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3228_o = n2905_o ? 1'b1 : n3227_o;
  assign n3229_o = enable_1[67];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3230_o = n2906_o ? 1'b1 : n3229_o;
  assign n3231_o = enable_1[68];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3232_o = n2907_o ? 1'b1 : n3231_o;
  assign n3233_o = enable_1[69];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3234_o = n2908_o ? 1'b1 : n3233_o;
  assign n3235_o = enable_1[70];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3236_o = n2909_o ? 1'b1 : n3235_o;
  assign n3237_o = enable_1[71];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3238_o = n2910_o ? 1'b1 : n3237_o;
  assign n3239_o = enable_1[72];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3240_o = n2911_o ? 1'b1 : n3239_o;
  assign n3241_o = enable_1[73];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3242_o = n2912_o ? 1'b1 : n3241_o;
  assign n3243_o = enable_1[74];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3244_o = n2913_o ? 1'b1 : n3243_o;
  assign n3245_o = enable_1[75];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3246_o = n2914_o ? 1'b1 : n3245_o;
  assign n3247_o = enable_1[76];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3248_o = n2915_o ? 1'b1 : n3247_o;
  assign n3249_o = enable_1[77];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3250_o = n2916_o ? 1'b1 : n3249_o;
  assign n3251_o = enable_1[78];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3252_o = n2917_o ? 1'b1 : n3251_o;
  assign n3253_o = enable_1[79];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3254_o = n2918_o ? 1'b1 : n3253_o;
  assign n3255_o = enable_1[80];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3256_o = n2919_o ? 1'b1 : n3255_o;
  assign n3257_o = enable_1[81];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3258_o = n2920_o ? 1'b1 : n3257_o;
  assign n3259_o = enable_1[82];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3260_o = n2921_o ? 1'b1 : n3259_o;
  assign n3261_o = enable_1[83];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3262_o = n2922_o ? 1'b1 : n3261_o;
  assign n3263_o = enable_1[84];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3264_o = n2923_o ? 1'b1 : n3263_o;
  assign n3265_o = enable_1[85];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3266_o = n2924_o ? 1'b1 : n3265_o;
  assign n3267_o = enable_1[86];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3268_o = n2925_o ? 1'b1 : n3267_o;
  assign n3269_o = enable_1[87];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3270_o = n2926_o ? 1'b1 : n3269_o;
  assign n3271_o = enable_1[88];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3272_o = n2927_o ? 1'b1 : n3271_o;
  assign n3273_o = enable_1[89];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3274_o = n2928_o ? 1'b1 : n3273_o;
  assign n3275_o = enable_1[90];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3276_o = n2929_o ? 1'b1 : n3275_o;
  assign n3277_o = enable_1[91];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3278_o = n2930_o ? 1'b1 : n3277_o;
  assign n3279_o = enable_1[92];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3280_o = n2931_o ? 1'b1 : n3279_o;
  assign n3281_o = enable_1[93];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3282_o = n2932_o ? 1'b1 : n3281_o;
  assign n3283_o = enable_1[94];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3284_o = n2933_o ? 1'b1 : n3283_o;
  assign n3285_o = enable_1[95];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3286_o = n2934_o ? 1'b1 : n3285_o;
  assign n3287_o = enable_1[96];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3288_o = n2935_o ? 1'b1 : n3287_o;
  assign n3289_o = enable_1[97];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3290_o = n2936_o ? 1'b1 : n3289_o;
  assign n3291_o = enable_1[98];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3292_o = n2937_o ? 1'b1 : n3291_o;
  assign n3293_o = enable_1[99];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3294_o = n2938_o ? 1'b1 : n3293_o;
  assign n3295_o = enable_1[100];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3296_o = n2939_o ? 1'b1 : n3295_o;
  assign n3297_o = enable_1[101];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3298_o = n2940_o ? 1'b1 : n3297_o;
  assign n3299_o = enable_1[102];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3300_o = n2941_o ? 1'b1 : n3299_o;
  assign n3301_o = enable_1[103];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3302_o = n2942_o ? 1'b1 : n3301_o;
  assign n3303_o = enable_1[104];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3304_o = n2943_o ? 1'b1 : n3303_o;
  assign n3305_o = enable_1[105];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3306_o = n2944_o ? 1'b1 : n3305_o;
  assign n3307_o = enable_1[106];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3308_o = n2945_o ? 1'b1 : n3307_o;
  assign n3309_o = enable_1[107];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3310_o = n2946_o ? 1'b1 : n3309_o;
  assign n3311_o = enable_1[108];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3312_o = n2947_o ? 1'b1 : n3311_o;
  assign n3313_o = enable_1[109];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3314_o = n2948_o ? 1'b1 : n3313_o;
  assign n3315_o = enable_1[110];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3316_o = n2949_o ? 1'b1 : n3315_o;
  assign n3317_o = enable_1[111];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3318_o = n2950_o ? 1'b1 : n3317_o;
  assign n3319_o = enable_1[112];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3320_o = n2951_o ? 1'b1 : n3319_o;
  assign n3321_o = enable_1[113];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3322_o = n2952_o ? 1'b1 : n3321_o;
  assign n3323_o = enable_1[114];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3324_o = n2953_o ? 1'b1 : n3323_o;
  assign n3325_o = enable_1[115];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3326_o = n2954_o ? 1'b1 : n3325_o;
  assign n3327_o = enable_1[116];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3328_o = n2955_o ? 1'b1 : n3327_o;
  assign n3329_o = enable_1[117];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3330_o = n2956_o ? 1'b1 : n3329_o;
  assign n3331_o = enable_1[118];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3332_o = n2957_o ? 1'b1 : n3331_o;
  assign n3333_o = enable_1[119];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3334_o = n2958_o ? 1'b1 : n3333_o;
  assign n3335_o = enable_1[120];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3336_o = n2959_o ? 1'b1 : n3335_o;
  assign n3337_o = enable_1[121];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3338_o = n2960_o ? 1'b1 : n3337_o;
  assign n3339_o = enable_1[122];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3340_o = n2961_o ? 1'b1 : n3339_o;
  assign n3341_o = enable_1[123];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3342_o = n2962_o ? 1'b1 : n3341_o;
  assign n3343_o = enable_1[124];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3344_o = n2963_o ? 1'b1 : n3343_o;
  assign n3345_o = enable_1[125];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3346_o = n2964_o ? 1'b1 : n3345_o;
  assign n3347_o = enable_1[126];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3348_o = n2965_o ? 1'b1 : n3347_o;
  assign n3349_o = enable_1[127];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3350_o = n2966_o ? 1'b1 : n3349_o;
  assign n3351_o = enable_1[128];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3352_o = n2967_o ? 1'b1 : n3351_o;
  assign n3353_o = enable_1[129];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3354_o = n2968_o ? 1'b1 : n3353_o;
  assign n3355_o = enable_1[130];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3356_o = n2969_o ? 1'b1 : n3355_o;
  assign n3357_o = enable_1[131];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3358_o = n2970_o ? 1'b1 : n3357_o;
  assign n3359_o = enable_1[132];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3360_o = n2971_o ? 1'b1 : n3359_o;
  assign n3361_o = enable_1[133];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3362_o = n2972_o ? 1'b1 : n3361_o;
  assign n3363_o = enable_1[134];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3364_o = n2973_o ? 1'b1 : n3363_o;
  assign n3365_o = enable_1[135];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3366_o = n2974_o ? 1'b1 : n3365_o;
  assign n3367_o = enable_1[136];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3368_o = n2975_o ? 1'b1 : n3367_o;
  assign n3369_o = enable_1[137];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3370_o = n2976_o ? 1'b1 : n3369_o;
  assign n3371_o = enable_1[138];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3372_o = n2977_o ? 1'b1 : n3371_o;
  assign n3373_o = enable_1[139];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3374_o = n2978_o ? 1'b1 : n3373_o;
  assign n3375_o = enable_1[140];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3376_o = n2979_o ? 1'b1 : n3375_o;
  assign n3377_o = enable_1[141];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3378_o = n2980_o ? 1'b1 : n3377_o;
  assign n3379_o = enable_1[142];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3380_o = n2981_o ? 1'b1 : n3379_o;
  assign n3381_o = enable_1[143];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3382_o = n2982_o ? 1'b1 : n3381_o;
  assign n3383_o = enable_1[144];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3384_o = n2983_o ? 1'b1 : n3383_o;
  assign n3385_o = enable_1[145];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3386_o = n2984_o ? 1'b1 : n3385_o;
  assign n3387_o = enable_1[146];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3388_o = n2985_o ? 1'b1 : n3387_o;
  assign n3389_o = enable_1[147];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3390_o = n2986_o ? 1'b1 : n3389_o;
  assign n3391_o = enable_1[148];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3392_o = n2987_o ? 1'b1 : n3391_o;
  assign n3393_o = enable_1[149];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3394_o = n2988_o ? 1'b1 : n3393_o;
  assign n3395_o = enable_1[150];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3396_o = n2989_o ? 1'b1 : n3395_o;
  assign n3397_o = enable_1[151];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3398_o = n2990_o ? 1'b1 : n3397_o;
  assign n3399_o = enable_1[152];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3400_o = n2991_o ? 1'b1 : n3399_o;
  assign n3401_o = enable_1[153];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3402_o = n2992_o ? 1'b1 : n3401_o;
  assign n3403_o = enable_1[154];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3404_o = n2993_o ? 1'b1 : n3403_o;
  assign n3405_o = enable_1[155];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3406_o = n2994_o ? 1'b1 : n3405_o;
  assign n3407_o = enable_1[156];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3408_o = n2995_o ? 1'b1 : n3407_o;
  assign n3409_o = enable_1[157];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3410_o = n2996_o ? 1'b1 : n3409_o;
  assign n3411_o = enable_1[158];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3412_o = n2997_o ? 1'b1 : n3411_o;
  assign n3413_o = enable_1[159];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3414_o = n2998_o ? 1'b1 : n3413_o;
  assign n3415_o = enable_1[160];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3416_o = n2999_o ? 1'b1 : n3415_o;
  assign n3417_o = enable_1[161];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3418_o = n3000_o ? 1'b1 : n3417_o;
  assign n3419_o = enable_1[162];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3420_o = n3001_o ? 1'b1 : n3419_o;
  assign n3421_o = enable_1[163];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3422_o = n3002_o ? 1'b1 : n3421_o;
  assign n3423_o = enable_1[164];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3424_o = n3003_o ? 1'b1 : n3423_o;
  assign n3425_o = enable_1[165];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3426_o = n3004_o ? 1'b1 : n3425_o;
  assign n3427_o = enable_1[166];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3428_o = n3005_o ? 1'b1 : n3427_o;
  assign n3429_o = enable_1[167];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3430_o = n3006_o ? 1'b1 : n3429_o;
  assign n3431_o = enable_1[168];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3432_o = n3007_o ? 1'b1 : n3431_o;
  assign n3433_o = enable_1[169];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3434_o = n3008_o ? 1'b1 : n3433_o;
  assign n3435_o = enable_1[170];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3436_o = n3009_o ? 1'b1 : n3435_o;
  assign n3437_o = enable_1[171];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3438_o = n3010_o ? 1'b1 : n3437_o;
  assign n3439_o = enable_1[172];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3440_o = n3011_o ? 1'b1 : n3439_o;
  assign n3441_o = enable_1[173];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3442_o = n3012_o ? 1'b1 : n3441_o;
  assign n3443_o = enable_1[174];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3444_o = n3013_o ? 1'b1 : n3443_o;
  assign n3445_o = enable_1[175];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3446_o = n3014_o ? 1'b1 : n3445_o;
  assign n3447_o = enable_1[176];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3448_o = n3015_o ? 1'b1 : n3447_o;
  assign n3449_o = enable_1[177];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3450_o = n3016_o ? 1'b1 : n3449_o;
  assign n3451_o = enable_1[178];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3452_o = n3017_o ? 1'b1 : n3451_o;
  assign n3453_o = enable_1[179];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3454_o = n3018_o ? 1'b1 : n3453_o;
  assign n3455_o = enable_1[180];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3456_o = n3019_o ? 1'b1 : n3455_o;
  assign n3457_o = enable_1[181];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3458_o = n3020_o ? 1'b1 : n3457_o;
  assign n3459_o = enable_1[182];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3460_o = n3021_o ? 1'b1 : n3459_o;
  assign n3461_o = enable_1[183];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3462_o = n3022_o ? 1'b1 : n3461_o;
  assign n3463_o = enable_1[184];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3464_o = n3023_o ? 1'b1 : n3463_o;
  assign n3465_o = enable_1[185];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3466_o = n3024_o ? 1'b1 : n3465_o;
  assign n3467_o = enable_1[186];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3468_o = n3025_o ? 1'b1 : n3467_o;
  assign n3469_o = enable_1[187];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3470_o = n3026_o ? 1'b1 : n3469_o;
  assign n3471_o = enable_1[188];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3472_o = n3027_o ? 1'b1 : n3471_o;
  assign n3473_o = enable_1[189];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3474_o = n3028_o ? 1'b1 : n3473_o;
  assign n3475_o = enable_1[190];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3476_o = n3029_o ? 1'b1 : n3475_o;
  assign n3477_o = enable_1[191];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3478_o = n3030_o ? 1'b1 : n3477_o;
  assign n3479_o = enable_1[192];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3480_o = n3031_o ? 1'b1 : n3479_o;
  assign n3481_o = enable_1[193];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3482_o = n3032_o ? 1'b1 : n3481_o;
  assign n3483_o = enable_1[194];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3484_o = n3033_o ? 1'b1 : n3483_o;
  assign n3485_o = enable_1[195];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3486_o = n3034_o ? 1'b1 : n3485_o;
  assign n3487_o = enable_1[196];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3488_o = n3035_o ? 1'b1 : n3487_o;
  assign n3489_o = enable_1[197];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3490_o = n3036_o ? 1'b1 : n3489_o;
  assign n3491_o = enable_1[198];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3492_o = n3037_o ? 1'b1 : n3491_o;
  assign n3493_o = enable_1[199];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3494_o = n3038_o ? 1'b1 : n3493_o;
  assign n3495_o = enable_1[200];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3496_o = n3039_o ? 1'b1 : n3495_o;
  assign n3497_o = enable_1[201];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3498_o = n3040_o ? 1'b1 : n3497_o;
  assign n3499_o = enable_1[202];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3500_o = n3041_o ? 1'b1 : n3499_o;
  assign n3501_o = enable_1[203];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3502_o = n3042_o ? 1'b1 : n3501_o;
  assign n3503_o = enable_1[204];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3504_o = n3043_o ? 1'b1 : n3503_o;
  assign n3505_o = enable_1[205];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3506_o = n3044_o ? 1'b1 : n3505_o;
  assign n3507_o = enable_1[206];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3508_o = n3045_o ? 1'b1 : n3507_o;
  assign n3509_o = enable_1[207];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3510_o = n3046_o ? 1'b1 : n3509_o;
  assign n3511_o = enable_1[208];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3512_o = n3047_o ? 1'b1 : n3511_o;
  assign n3513_o = enable_1[209];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3514_o = n3048_o ? 1'b1 : n3513_o;
  assign n3515_o = enable_1[210];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3516_o = n3049_o ? 1'b1 : n3515_o;
  assign n3517_o = enable_1[211];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3518_o = n3050_o ? 1'b1 : n3517_o;
  assign n3519_o = enable_1[212];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3520_o = n3051_o ? 1'b1 : n3519_o;
  assign n3521_o = enable_1[213];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3522_o = n3052_o ? 1'b1 : n3521_o;
  assign n3523_o = enable_1[214];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3524_o = n3053_o ? 1'b1 : n3523_o;
  assign n3525_o = enable_1[215];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3526_o = n3054_o ? 1'b1 : n3525_o;
  assign n3527_o = enable_1[216];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3528_o = n3055_o ? 1'b1 : n3527_o;
  assign n3529_o = enable_1[217];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3530_o = n3056_o ? 1'b1 : n3529_o;
  assign n3531_o = enable_1[218];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3532_o = n3057_o ? 1'b1 : n3531_o;
  assign n3533_o = enable_1[219];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3534_o = n3058_o ? 1'b1 : n3533_o;
  assign n3535_o = enable_1[220];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3536_o = n3059_o ? 1'b1 : n3535_o;
  assign n3537_o = enable_1[221];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3538_o = n3060_o ? 1'b1 : n3537_o;
  assign n3539_o = enable_1[222];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3540_o = n3061_o ? 1'b1 : n3539_o;
  assign n3541_o = enable_1[223];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3542_o = n3062_o ? 1'b1 : n3541_o;
  assign n3543_o = enable_1[224];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3544_o = n3063_o ? 1'b1 : n3543_o;
  assign n3545_o = enable_1[225];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3546_o = n3064_o ? 1'b1 : n3545_o;
  assign n3547_o = enable_1[226];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3548_o = n3065_o ? 1'b1 : n3547_o;
  assign n3549_o = enable_1[227];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3550_o = n3066_o ? 1'b1 : n3549_o;
  assign n3551_o = enable_1[228];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3552_o = n3067_o ? 1'b1 : n3551_o;
  assign n3553_o = enable_1[229];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3554_o = n3068_o ? 1'b1 : n3553_o;
  assign n3555_o = enable_1[230];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3556_o = n3069_o ? 1'b1 : n3555_o;
  assign n3557_o = enable_1[231];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3558_o = n3070_o ? 1'b1 : n3557_o;
  assign n3559_o = enable_1[232];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3560_o = n3071_o ? 1'b1 : n3559_o;
  assign n3561_o = enable_1[233];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3562_o = n3072_o ? 1'b1 : n3561_o;
  assign n3563_o = enable_1[234];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3564_o = n3073_o ? 1'b1 : n3563_o;
  assign n3565_o = enable_1[235];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3566_o = n3074_o ? 1'b1 : n3565_o;
  assign n3567_o = enable_1[236];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3568_o = n3075_o ? 1'b1 : n3567_o;
  assign n3569_o = enable_1[237];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3570_o = n3076_o ? 1'b1 : n3569_o;
  assign n3571_o = enable_1[238];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3572_o = n3077_o ? 1'b1 : n3571_o;
  assign n3573_o = enable_1[239];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3574_o = n3078_o ? 1'b1 : n3573_o;
  assign n3575_o = enable_1[240];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3576_o = n3079_o ? 1'b1 : n3575_o;
  assign n3577_o = enable_1[241];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3578_o = n3080_o ? 1'b1 : n3577_o;
  assign n3579_o = enable_1[242];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3580_o = n3081_o ? 1'b1 : n3579_o;
  assign n3581_o = enable_1[243];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3582_o = n3082_o ? 1'b1 : n3581_o;
  assign n3583_o = enable_1[244];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3584_o = n3083_o ? 1'b1 : n3583_o;
  assign n3585_o = enable_1[245];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3586_o = n3084_o ? 1'b1 : n3585_o;
  assign n3587_o = enable_1[246];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3588_o = n3085_o ? 1'b1 : n3587_o;
  assign n3589_o = enable_1[247];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3590_o = n3086_o ? 1'b1 : n3589_o;
  assign n3591_o = enable_1[248];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3592_o = n3087_o ? 1'b1 : n3591_o;
  assign n3593_o = enable_1[249];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3594_o = n3088_o ? 1'b1 : n3593_o;
  assign n3595_o = enable_1[250];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3596_o = n3089_o ? 1'b1 : n3595_o;
  assign n3597_o = enable_1[251];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3598_o = n3090_o ? 1'b1 : n3597_o;
  assign n3599_o = enable_1[252];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3600_o = n3091_o ? 1'b1 : n3599_o;
  assign n3601_o = enable_1[253];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3602_o = n3092_o ? 1'b1 : n3601_o;
  assign n3603_o = enable_1[254];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3604_o = n3093_o ? 1'b1 : n3603_o;
  assign n3605_o = enable_1[255];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:437:21  */
  assign n3606_o = n3094_o ? 1'b1 : n3605_o;
  assign n3607_o = {n3606_o, n3604_o, n3602_o, n3600_o, n3598_o, n3596_o, n3594_o, n3592_o, n3590_o, n3588_o, n3586_o, n3584_o, n3582_o, n3580_o, n3578_o, n3576_o, n3574_o, n3572_o, n3570_o, n3568_o, n3566_o, n3564_o, n3562_o, n3560_o, n3558_o, n3556_o, n3554_o, n3552_o, n3550_o, n3548_o, n3546_o, n3544_o, n3542_o, n3540_o, n3538_o, n3536_o, n3534_o, n3532_o, n3530_o, n3528_o, n3526_o, n3524_o, n3522_o, n3520_o, n3518_o, n3516_o, n3514_o, n3512_o, n3510_o, n3508_o, n3506_o, n3504_o, n3502_o, n3500_o, n3498_o, n3496_o, n3494_o, n3492_o, n3490_o, n3488_o, n3486_o, n3484_o, n3482_o, n3480_o, n3478_o, n3476_o, n3474_o, n3472_o, n3470_o, n3468_o, n3466_o, n3464_o, n3462_o, n3460_o, n3458_o, n3456_o, n3454_o, n3452_o, n3450_o, n3448_o, n3446_o, n3444_o, n3442_o, n3440_o, n3438_o, n3436_o, n3434_o, n3432_o, n3430_o, n3428_o, n3426_o, n3424_o, n3422_o, n3420_o, n3418_o, n3416_o, n3414_o, n3412_o, n3410_o, n3408_o, n3406_o, n3404_o, n3402_o, n3400_o, n3398_o, n3396_o, n3394_o, n3392_o, n3390_o, n3388_o, n3386_o, n3384_o, n3382_o, n3380_o, n3378_o, n3376_o, n3374_o, n3372_o, n3370_o, n3368_o, n3366_o, n3364_o, n3362_o, n3360_o, n3358_o, n3356_o, n3354_o, n3352_o, n3350_o, n3348_o, n3346_o, n3344_o, n3342_o, n3340_o, n3338_o, n3336_o, n3334_o, n3332_o, n3330_o, n3328_o, n3326_o, n3324_o, n3322_o, n3320_o, n3318_o, n3316_o, n3314_o, n3312_o, n3310_o, n3308_o, n3306_o, n3304_o, n3302_o, n3300_o, n3298_o, n3296_o, n3294_o, n3292_o, n3290_o, n3288_o, n3286_o, n3284_o, n3282_o, n3280_o, n3278_o, n3276_o, n3274_o, n3272_o, n3270_o, n3268_o, n3266_o, n3264_o, n3262_o, n3260_o, n3258_o, n3256_o, n3254_o, n3252_o, n3250_o, n3248_o, n3246_o, n3244_o, n3242_o, n3240_o, n3238_o, n3236_o, n3234_o, n3232_o, n3230_o, n3228_o, n3226_o, n3224_o, n3222_o, n3220_o, n3218_o, n3216_o, n3214_o, n3212_o, n3210_o, n3208_o, n3206_o, n3204_o, n3202_o, n3200_o, n3198_o, n3196_o, n3194_o, n3192_o, n3190_o, n3188_o, n3186_o, n3184_o, n3182_o, n3180_o, n3178_o, n3176_o, n3174_o, n3172_o, n3170_o, n3168_o, n3166_o, n3164_o, n3162_o, n3160_o, n3158_o, n3156_o, n3154_o, n3152_o, n3150_o, n3148_o, n3146_o, n3144_o, n3142_o, n3140_o, n3138_o, n3136_o, n3134_o, n3132_o, n3130_o, n3128_o, n3126_o, n3124_o, n3122_o, n3120_o, n3118_o, n3116_o, n3114_o, n3112_o, n3110_o, n3108_o, n3106_o, n3104_o, n3102_o, n3100_o, n3098_o, n3096_o};
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3608_o = n267_o[7];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3609_o = ~n3608_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3610_o = n267_o[6];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3611_o = ~n3610_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3612_o = n3609_o & n3611_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3613_o = n3609_o & n3610_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3614_o = n3608_o & n3611_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3615_o = n3608_o & n3610_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3616_o = n267_o[5];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3617_o = ~n3616_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3618_o = n3612_o & n3617_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3619_o = n3612_o & n3616_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3620_o = n3613_o & n3617_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3621_o = n3613_o & n3616_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3622_o = n3614_o & n3617_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3623_o = n3614_o & n3616_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3624_o = n3615_o & n3617_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3625_o = n3615_o & n3616_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3626_o = n267_o[4];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3627_o = ~n3626_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3628_o = n3618_o & n3627_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3629_o = n3618_o & n3626_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3630_o = n3619_o & n3627_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3631_o = n3619_o & n3626_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3632_o = n3620_o & n3627_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3633_o = n3620_o & n3626_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3634_o = n3621_o & n3627_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3635_o = n3621_o & n3626_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3636_o = n3622_o & n3627_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3637_o = n3622_o & n3626_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3638_o = n3623_o & n3627_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3639_o = n3623_o & n3626_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3640_o = n3624_o & n3627_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3641_o = n3624_o & n3626_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3642_o = n3625_o & n3627_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3643_o = n3625_o & n3626_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3644_o = n267_o[3];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3645_o = ~n3644_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3646_o = n3628_o & n3645_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3647_o = n3628_o & n3644_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3648_o = n3629_o & n3645_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3649_o = n3629_o & n3644_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3650_o = n3630_o & n3645_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3651_o = n3630_o & n3644_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3652_o = n3631_o & n3645_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3653_o = n3631_o & n3644_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3654_o = n3632_o & n3645_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3655_o = n3632_o & n3644_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3656_o = n3633_o & n3645_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3657_o = n3633_o & n3644_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3658_o = n3634_o & n3645_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3659_o = n3634_o & n3644_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3660_o = n3635_o & n3645_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3661_o = n3635_o & n3644_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3662_o = n3636_o & n3645_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3663_o = n3636_o & n3644_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3664_o = n3637_o & n3645_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3665_o = n3637_o & n3644_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3666_o = n3638_o & n3645_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3667_o = n3638_o & n3644_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3668_o = n3639_o & n3645_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3669_o = n3639_o & n3644_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3670_o = n3640_o & n3645_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3671_o = n3640_o & n3644_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3672_o = n3641_o & n3645_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3673_o = n3641_o & n3644_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3674_o = n3642_o & n3645_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3675_o = n3642_o & n3644_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3676_o = n3643_o & n3645_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3677_o = n3643_o & n3644_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3678_o = n267_o[2];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3679_o = ~n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3680_o = n3646_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3681_o = n3646_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3682_o = n3647_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3683_o = n3647_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3684_o = n3648_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3685_o = n3648_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3686_o = n3649_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3687_o = n3649_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3688_o = n3650_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3689_o = n3650_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3690_o = n3651_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3691_o = n3651_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3692_o = n3652_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3693_o = n3652_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3694_o = n3653_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3695_o = n3653_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3696_o = n3654_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3697_o = n3654_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3698_o = n3655_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3699_o = n3655_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3700_o = n3656_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3701_o = n3656_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3702_o = n3657_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3703_o = n3657_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3704_o = n3658_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3705_o = n3658_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3706_o = n3659_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3707_o = n3659_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3708_o = n3660_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3709_o = n3660_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3710_o = n3661_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3711_o = n3661_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3712_o = n3662_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3713_o = n3662_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3714_o = n3663_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3715_o = n3663_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3716_o = n3664_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3717_o = n3664_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3718_o = n3665_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3719_o = n3665_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3720_o = n3666_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3721_o = n3666_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3722_o = n3667_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3723_o = n3667_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3724_o = n3668_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3725_o = n3668_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3726_o = n3669_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3727_o = n3669_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3728_o = n3670_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3729_o = n3670_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3730_o = n3671_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3731_o = n3671_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3732_o = n3672_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3733_o = n3672_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3734_o = n3673_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3735_o = n3673_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3736_o = n3674_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3737_o = n3674_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3738_o = n3675_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3739_o = n3675_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3740_o = n3676_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3741_o = n3676_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3742_o = n3677_o & n3679_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3743_o = n3677_o & n3678_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3744_o = n267_o[1];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3745_o = ~n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3746_o = n3680_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3747_o = n3680_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3748_o = n3681_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3749_o = n3681_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3750_o = n3682_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3751_o = n3682_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3752_o = n3683_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3753_o = n3683_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3754_o = n3684_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3755_o = n3684_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3756_o = n3685_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3757_o = n3685_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3758_o = n3686_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3759_o = n3686_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3760_o = n3687_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3761_o = n3687_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3762_o = n3688_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3763_o = n3688_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3764_o = n3689_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3765_o = n3689_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3766_o = n3690_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3767_o = n3690_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3768_o = n3691_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3769_o = n3691_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3770_o = n3692_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3771_o = n3692_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3772_o = n3693_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3773_o = n3693_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3774_o = n3694_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3775_o = n3694_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3776_o = n3695_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3777_o = n3695_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3778_o = n3696_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3779_o = n3696_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3780_o = n3697_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3781_o = n3697_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3782_o = n3698_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3783_o = n3698_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3784_o = n3699_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3785_o = n3699_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3786_o = n3700_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3787_o = n3700_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3788_o = n3701_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3789_o = n3701_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3790_o = n3702_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3791_o = n3702_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3792_o = n3703_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3793_o = n3703_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3794_o = n3704_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3795_o = n3704_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3796_o = n3705_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3797_o = n3705_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3798_o = n3706_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3799_o = n3706_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3800_o = n3707_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3801_o = n3707_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3802_o = n3708_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3803_o = n3708_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3804_o = n3709_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3805_o = n3709_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3806_o = n3710_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3807_o = n3710_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3808_o = n3711_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3809_o = n3711_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3810_o = n3712_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3811_o = n3712_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3812_o = n3713_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3813_o = n3713_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3814_o = n3714_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3815_o = n3714_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3816_o = n3715_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3817_o = n3715_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3818_o = n3716_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3819_o = n3716_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3820_o = n3717_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3821_o = n3717_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3822_o = n3718_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3823_o = n3718_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3824_o = n3719_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3825_o = n3719_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3826_o = n3720_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3827_o = n3720_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3828_o = n3721_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3829_o = n3721_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3830_o = n3722_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3831_o = n3722_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3832_o = n3723_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3833_o = n3723_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3834_o = n3724_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3835_o = n3724_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3836_o = n3725_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3837_o = n3725_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3838_o = n3726_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3839_o = n3726_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3840_o = n3727_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3841_o = n3727_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3842_o = n3728_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3843_o = n3728_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3844_o = n3729_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3845_o = n3729_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3846_o = n3730_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3847_o = n3730_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3848_o = n3731_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3849_o = n3731_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3850_o = n3732_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3851_o = n3732_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3852_o = n3733_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3853_o = n3733_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3854_o = n3734_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3855_o = n3734_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3856_o = n3735_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3857_o = n3735_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3858_o = n3736_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3859_o = n3736_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3860_o = n3737_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3861_o = n3737_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3862_o = n3738_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3863_o = n3738_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3864_o = n3739_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3865_o = n3739_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3866_o = n3740_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3867_o = n3740_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3868_o = n3741_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3869_o = n3741_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3870_o = n3742_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3871_o = n3742_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3872_o = n3743_o & n3745_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3873_o = n3743_o & n3744_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3874_o = n267_o[0];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3875_o = ~n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3876_o = n3746_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3877_o = n3746_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3878_o = n3747_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3879_o = n3747_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3880_o = n3748_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3881_o = n3748_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3882_o = n3749_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3883_o = n3749_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3884_o = n3750_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3885_o = n3750_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3886_o = n3751_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3887_o = n3751_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3888_o = n3752_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3889_o = n3752_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3890_o = n3753_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3891_o = n3753_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3892_o = n3754_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3893_o = n3754_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3894_o = n3755_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3895_o = n3755_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3896_o = n3756_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3897_o = n3756_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3898_o = n3757_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3899_o = n3757_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3900_o = n3758_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3901_o = n3758_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3902_o = n3759_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3903_o = n3759_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3904_o = n3760_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3905_o = n3760_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3906_o = n3761_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3907_o = n3761_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3908_o = n3762_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3909_o = n3762_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3910_o = n3763_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3911_o = n3763_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3912_o = n3764_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3913_o = n3764_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3914_o = n3765_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3915_o = n3765_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3916_o = n3766_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3917_o = n3766_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3918_o = n3767_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3919_o = n3767_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3920_o = n3768_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3921_o = n3768_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3922_o = n3769_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3923_o = n3769_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3924_o = n3770_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3925_o = n3770_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3926_o = n3771_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3927_o = n3771_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3928_o = n3772_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3929_o = n3772_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3930_o = n3773_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3931_o = n3773_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3932_o = n3774_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3933_o = n3774_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3934_o = n3775_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3935_o = n3775_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3936_o = n3776_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3937_o = n3776_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3938_o = n3777_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3939_o = n3777_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3940_o = n3778_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3941_o = n3778_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3942_o = n3779_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3943_o = n3779_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3944_o = n3780_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3945_o = n3780_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3946_o = n3781_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3947_o = n3781_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3948_o = n3782_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3949_o = n3782_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3950_o = n3783_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3951_o = n3783_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3952_o = n3784_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3953_o = n3784_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3954_o = n3785_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3955_o = n3785_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3956_o = n3786_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3957_o = n3786_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3958_o = n3787_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3959_o = n3787_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3960_o = n3788_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3961_o = n3788_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3962_o = n3789_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3963_o = n3789_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3964_o = n3790_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3965_o = n3790_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3966_o = n3791_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3967_o = n3791_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3968_o = n3792_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3969_o = n3792_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3970_o = n3793_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3971_o = n3793_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3972_o = n3794_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3973_o = n3794_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3974_o = n3795_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3975_o = n3795_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3976_o = n3796_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3977_o = n3796_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3978_o = n3797_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3979_o = n3797_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3980_o = n3798_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3981_o = n3798_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3982_o = n3799_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3983_o = n3799_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3984_o = n3800_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3985_o = n3800_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3986_o = n3801_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3987_o = n3801_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3988_o = n3802_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3989_o = n3802_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3990_o = n3803_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3991_o = n3803_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3992_o = n3804_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3993_o = n3804_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3994_o = n3805_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3995_o = n3805_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3996_o = n3806_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3997_o = n3806_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3998_o = n3807_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n3999_o = n3807_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4000_o = n3808_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4001_o = n3808_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4002_o = n3809_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4003_o = n3809_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4004_o = n3810_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4005_o = n3810_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4006_o = n3811_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4007_o = n3811_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4008_o = n3812_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4009_o = n3812_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4010_o = n3813_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4011_o = n3813_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4012_o = n3814_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4013_o = n3814_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4014_o = n3815_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4015_o = n3815_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4016_o = n3816_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4017_o = n3816_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4018_o = n3817_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4019_o = n3817_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4020_o = n3818_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4021_o = n3818_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4022_o = n3819_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4023_o = n3819_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4024_o = n3820_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4025_o = n3820_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4026_o = n3821_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4027_o = n3821_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4028_o = n3822_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4029_o = n3822_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4030_o = n3823_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4031_o = n3823_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4032_o = n3824_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4033_o = n3824_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4034_o = n3825_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4035_o = n3825_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4036_o = n3826_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4037_o = n3826_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4038_o = n3827_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4039_o = n3827_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4040_o = n3828_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4041_o = n3828_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4042_o = n3829_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4043_o = n3829_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4044_o = n3830_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4045_o = n3830_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4046_o = n3831_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4047_o = n3831_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4048_o = n3832_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4049_o = n3832_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4050_o = n3833_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4051_o = n3833_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4052_o = n3834_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4053_o = n3834_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4054_o = n3835_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4055_o = n3835_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4056_o = n3836_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4057_o = n3836_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4058_o = n3837_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4059_o = n3837_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4060_o = n3838_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4061_o = n3838_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4062_o = n3839_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4063_o = n3839_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4064_o = n3840_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4065_o = n3840_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4066_o = n3841_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4067_o = n3841_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4068_o = n3842_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4069_o = n3842_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4070_o = n3843_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4071_o = n3843_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4072_o = n3844_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4073_o = n3844_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4074_o = n3845_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4075_o = n3845_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4076_o = n3846_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4077_o = n3846_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4078_o = n3847_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4079_o = n3847_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4080_o = n3848_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4081_o = n3848_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4082_o = n3849_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4083_o = n3849_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4084_o = n3850_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4085_o = n3850_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4086_o = n3851_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4087_o = n3851_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4088_o = n3852_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4089_o = n3852_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4090_o = n3853_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4091_o = n3853_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4092_o = n3854_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4093_o = n3854_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4094_o = n3855_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4095_o = n3855_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4096_o = n3856_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4097_o = n3856_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4098_o = n3857_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4099_o = n3857_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4100_o = n3858_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4101_o = n3858_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4102_o = n3859_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4103_o = n3859_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4104_o = n3860_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4105_o = n3860_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4106_o = n3861_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4107_o = n3861_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4108_o = n3862_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4109_o = n3862_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4110_o = n3863_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4111_o = n3863_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4112_o = n3864_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4113_o = n3864_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4114_o = n3865_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4115_o = n3865_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4116_o = n3866_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4117_o = n3866_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4118_o = n3867_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4119_o = n3867_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4120_o = n3868_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4121_o = n3868_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4122_o = n3869_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4123_o = n3869_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4124_o = n3870_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4125_o = n3870_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4126_o = n3871_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4127_o = n3871_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4128_o = n3872_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4129_o = n3872_o & n3874_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4130_o = n3873_o & n3875_o;
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4131_o = n3873_o & n3874_o;
  assign n4132_o = enable_2[0];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4133_o = n3876_o ? 1'b1 : n4132_o;
  assign n4134_o = enable_2[1];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4135_o = n3877_o ? 1'b1 : n4134_o;
  assign n4136_o = enable_2[2];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4137_o = n3878_o ? 1'b1 : n4136_o;
  assign n4138_o = enable_2[3];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4139_o = n3879_o ? 1'b1 : n4138_o;
  assign n4140_o = enable_2[4];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4141_o = n3880_o ? 1'b1 : n4140_o;
  assign n4142_o = enable_2[5];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4143_o = n3881_o ? 1'b1 : n4142_o;
  assign n4144_o = enable_2[6];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4145_o = n3882_o ? 1'b1 : n4144_o;
  assign n4146_o = enable_2[7];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4147_o = n3883_o ? 1'b1 : n4146_o;
  assign n4148_o = enable_2[8];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4149_o = n3884_o ? 1'b1 : n4148_o;
  assign n4150_o = enable_2[9];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4151_o = n3885_o ? 1'b1 : n4150_o;
  assign n4152_o = enable_2[10];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4153_o = n3886_o ? 1'b1 : n4152_o;
  assign n4154_o = enable_2[11];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4155_o = n3887_o ? 1'b1 : n4154_o;
  assign n4156_o = enable_2[12];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4157_o = n3888_o ? 1'b1 : n4156_o;
  assign n4158_o = enable_2[13];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4159_o = n3889_o ? 1'b1 : n4158_o;
  assign n4160_o = enable_2[14];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4161_o = n3890_o ? 1'b1 : n4160_o;
  assign n4162_o = enable_2[15];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4163_o = n3891_o ? 1'b1 : n4162_o;
  assign n4164_o = enable_2[16];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4165_o = n3892_o ? 1'b1 : n4164_o;
  assign n4166_o = enable_2[17];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4167_o = n3893_o ? 1'b1 : n4166_o;
  assign n4168_o = enable_2[18];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4169_o = n3894_o ? 1'b1 : n4168_o;
  assign n4170_o = enable_2[19];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4171_o = n3895_o ? 1'b1 : n4170_o;
  assign n4172_o = enable_2[20];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4173_o = n3896_o ? 1'b1 : n4172_o;
  assign n4174_o = enable_2[21];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4175_o = n3897_o ? 1'b1 : n4174_o;
  assign n4176_o = enable_2[22];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4177_o = n3898_o ? 1'b1 : n4176_o;
  assign n4178_o = enable_2[23];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4179_o = n3899_o ? 1'b1 : n4178_o;
  assign n4180_o = enable_2[24];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4181_o = n3900_o ? 1'b1 : n4180_o;
  assign n4182_o = enable_2[25];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4183_o = n3901_o ? 1'b1 : n4182_o;
  assign n4184_o = enable_2[26];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4185_o = n3902_o ? 1'b1 : n4184_o;
  assign n4186_o = enable_2[27];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4187_o = n3903_o ? 1'b1 : n4186_o;
  assign n4188_o = enable_2[28];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4189_o = n3904_o ? 1'b1 : n4188_o;
  assign n4190_o = enable_2[29];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4191_o = n3905_o ? 1'b1 : n4190_o;
  assign n4192_o = enable_2[30];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4193_o = n3906_o ? 1'b1 : n4192_o;
  assign n4194_o = enable_2[31];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4195_o = n3907_o ? 1'b1 : n4194_o;
  assign n4196_o = enable_2[32];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4197_o = n3908_o ? 1'b1 : n4196_o;
  assign n4198_o = enable_2[33];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4199_o = n3909_o ? 1'b1 : n4198_o;
  assign n4200_o = enable_2[34];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4201_o = n3910_o ? 1'b1 : n4200_o;
  assign n4202_o = enable_2[35];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4203_o = n3911_o ? 1'b1 : n4202_o;
  assign n4204_o = enable_2[36];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4205_o = n3912_o ? 1'b1 : n4204_o;
  assign n4206_o = enable_2[37];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4207_o = n3913_o ? 1'b1 : n4206_o;
  assign n4208_o = enable_2[38];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4209_o = n3914_o ? 1'b1 : n4208_o;
  assign n4210_o = enable_2[39];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4211_o = n3915_o ? 1'b1 : n4210_o;
  assign n4212_o = enable_2[40];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4213_o = n3916_o ? 1'b1 : n4212_o;
  assign n4214_o = enable_2[41];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4215_o = n3917_o ? 1'b1 : n4214_o;
  assign n4216_o = enable_2[42];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4217_o = n3918_o ? 1'b1 : n4216_o;
  assign n4218_o = enable_2[43];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4219_o = n3919_o ? 1'b1 : n4218_o;
  assign n4220_o = enable_2[44];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4221_o = n3920_o ? 1'b1 : n4220_o;
  assign n4222_o = enable_2[45];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4223_o = n3921_o ? 1'b1 : n4222_o;
  assign n4224_o = enable_2[46];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4225_o = n3922_o ? 1'b1 : n4224_o;
  assign n4226_o = enable_2[47];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4227_o = n3923_o ? 1'b1 : n4226_o;
  assign n4228_o = enable_2[48];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4229_o = n3924_o ? 1'b1 : n4228_o;
  assign n4230_o = enable_2[49];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4231_o = n3925_o ? 1'b1 : n4230_o;
  assign n4232_o = enable_2[50];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4233_o = n3926_o ? 1'b1 : n4232_o;
  assign n4234_o = enable_2[51];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4235_o = n3927_o ? 1'b1 : n4234_o;
  assign n4236_o = enable_2[52];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4237_o = n3928_o ? 1'b1 : n4236_o;
  assign n4238_o = enable_2[53];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4239_o = n3929_o ? 1'b1 : n4238_o;
  assign n4240_o = enable_2[54];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4241_o = n3930_o ? 1'b1 : n4240_o;
  assign n4242_o = enable_2[55];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4243_o = n3931_o ? 1'b1 : n4242_o;
  assign n4244_o = enable_2[56];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4245_o = n3932_o ? 1'b1 : n4244_o;
  assign n4246_o = enable_2[57];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4247_o = n3933_o ? 1'b1 : n4246_o;
  assign n4248_o = enable_2[58];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4249_o = n3934_o ? 1'b1 : n4248_o;
  assign n4250_o = enable_2[59];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4251_o = n3935_o ? 1'b1 : n4250_o;
  assign n4252_o = enable_2[60];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4253_o = n3936_o ? 1'b1 : n4252_o;
  assign n4254_o = enable_2[61];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4255_o = n3937_o ? 1'b1 : n4254_o;
  assign n4256_o = enable_2[62];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4257_o = n3938_o ? 1'b1 : n4256_o;
  assign n4258_o = enable_2[63];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4259_o = n3939_o ? 1'b1 : n4258_o;
  assign n4260_o = enable_2[64];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4261_o = n3940_o ? 1'b1 : n4260_o;
  assign n4262_o = enable_2[65];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4263_o = n3941_o ? 1'b1 : n4262_o;
  assign n4264_o = enable_2[66];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4265_o = n3942_o ? 1'b1 : n4264_o;
  assign n4266_o = enable_2[67];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4267_o = n3943_o ? 1'b1 : n4266_o;
  assign n4268_o = enable_2[68];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4269_o = n3944_o ? 1'b1 : n4268_o;
  assign n4270_o = enable_2[69];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4271_o = n3945_o ? 1'b1 : n4270_o;
  assign n4272_o = enable_2[70];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4273_o = n3946_o ? 1'b1 : n4272_o;
  assign n4274_o = enable_2[71];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4275_o = n3947_o ? 1'b1 : n4274_o;
  assign n4276_o = enable_2[72];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4277_o = n3948_o ? 1'b1 : n4276_o;
  assign n4278_o = enable_2[73];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4279_o = n3949_o ? 1'b1 : n4278_o;
  assign n4280_o = enable_2[74];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4281_o = n3950_o ? 1'b1 : n4280_o;
  assign n4282_o = enable_2[75];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4283_o = n3951_o ? 1'b1 : n4282_o;
  assign n4284_o = enable_2[76];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4285_o = n3952_o ? 1'b1 : n4284_o;
  assign n4286_o = enable_2[77];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4287_o = n3953_o ? 1'b1 : n4286_o;
  assign n4288_o = enable_2[78];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4289_o = n3954_o ? 1'b1 : n4288_o;
  assign n4290_o = enable_2[79];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4291_o = n3955_o ? 1'b1 : n4290_o;
  assign n4292_o = enable_2[80];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4293_o = n3956_o ? 1'b1 : n4292_o;
  assign n4294_o = enable_2[81];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4295_o = n3957_o ? 1'b1 : n4294_o;
  assign n4296_o = enable_2[82];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4297_o = n3958_o ? 1'b1 : n4296_o;
  assign n4298_o = enable_2[83];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4299_o = n3959_o ? 1'b1 : n4298_o;
  assign n4300_o = enable_2[84];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4301_o = n3960_o ? 1'b1 : n4300_o;
  assign n4302_o = enable_2[85];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4303_o = n3961_o ? 1'b1 : n4302_o;
  assign n4304_o = enable_2[86];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4305_o = n3962_o ? 1'b1 : n4304_o;
  assign n4306_o = enable_2[87];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4307_o = n3963_o ? 1'b1 : n4306_o;
  assign n4308_o = enable_2[88];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4309_o = n3964_o ? 1'b1 : n4308_o;
  assign n4310_o = enable_2[89];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4311_o = n3965_o ? 1'b1 : n4310_o;
  assign n4312_o = enable_2[90];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4313_o = n3966_o ? 1'b1 : n4312_o;
  assign n4314_o = enable_2[91];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4315_o = n3967_o ? 1'b1 : n4314_o;
  assign n4316_o = enable_2[92];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4317_o = n3968_o ? 1'b1 : n4316_o;
  assign n4318_o = enable_2[93];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4319_o = n3969_o ? 1'b1 : n4318_o;
  assign n4320_o = enable_2[94];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4321_o = n3970_o ? 1'b1 : n4320_o;
  assign n4322_o = enable_2[95];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4323_o = n3971_o ? 1'b1 : n4322_o;
  assign n4324_o = enable_2[96];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4325_o = n3972_o ? 1'b1 : n4324_o;
  assign n4326_o = enable_2[97];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4327_o = n3973_o ? 1'b1 : n4326_o;
  assign n4328_o = enable_2[98];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4329_o = n3974_o ? 1'b1 : n4328_o;
  assign n4330_o = enable_2[99];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4331_o = n3975_o ? 1'b1 : n4330_o;
  assign n4332_o = enable_2[100];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4333_o = n3976_o ? 1'b1 : n4332_o;
  assign n4334_o = enable_2[101];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4335_o = n3977_o ? 1'b1 : n4334_o;
  assign n4336_o = enable_2[102];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4337_o = n3978_o ? 1'b1 : n4336_o;
  assign n4338_o = enable_2[103];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4339_o = n3979_o ? 1'b1 : n4338_o;
  assign n4340_o = enable_2[104];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4341_o = n3980_o ? 1'b1 : n4340_o;
  assign n4342_o = enable_2[105];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4343_o = n3981_o ? 1'b1 : n4342_o;
  assign n4344_o = enable_2[106];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4345_o = n3982_o ? 1'b1 : n4344_o;
  assign n4346_o = enable_2[107];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4347_o = n3983_o ? 1'b1 : n4346_o;
  assign n4348_o = enable_2[108];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4349_o = n3984_o ? 1'b1 : n4348_o;
  assign n4350_o = enable_2[109];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4351_o = n3985_o ? 1'b1 : n4350_o;
  assign n4352_o = enable_2[110];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4353_o = n3986_o ? 1'b1 : n4352_o;
  assign n4354_o = enable_2[111];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4355_o = n3987_o ? 1'b1 : n4354_o;
  assign n4356_o = enable_2[112];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4357_o = n3988_o ? 1'b1 : n4356_o;
  assign n4358_o = enable_2[113];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4359_o = n3989_o ? 1'b1 : n4358_o;
  assign n4360_o = enable_2[114];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4361_o = n3990_o ? 1'b1 : n4360_o;
  assign n4362_o = enable_2[115];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4363_o = n3991_o ? 1'b1 : n4362_o;
  assign n4364_o = enable_2[116];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4365_o = n3992_o ? 1'b1 : n4364_o;
  assign n4366_o = enable_2[117];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4367_o = n3993_o ? 1'b1 : n4366_o;
  assign n4368_o = enable_2[118];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4369_o = n3994_o ? 1'b1 : n4368_o;
  assign n4370_o = enable_2[119];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4371_o = n3995_o ? 1'b1 : n4370_o;
  assign n4372_o = enable_2[120];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4373_o = n3996_o ? 1'b1 : n4372_o;
  assign n4374_o = enable_2[121];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4375_o = n3997_o ? 1'b1 : n4374_o;
  assign n4376_o = enable_2[122];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4377_o = n3998_o ? 1'b1 : n4376_o;
  assign n4378_o = enable_2[123];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4379_o = n3999_o ? 1'b1 : n4378_o;
  assign n4380_o = enable_2[124];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4381_o = n4000_o ? 1'b1 : n4380_o;
  assign n4382_o = enable_2[125];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4383_o = n4001_o ? 1'b1 : n4382_o;
  assign n4384_o = enable_2[126];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4385_o = n4002_o ? 1'b1 : n4384_o;
  assign n4386_o = enable_2[127];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4387_o = n4003_o ? 1'b1 : n4386_o;
  assign n4388_o = enable_2[128];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4389_o = n4004_o ? 1'b1 : n4388_o;
  assign n4390_o = enable_2[129];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4391_o = n4005_o ? 1'b1 : n4390_o;
  assign n4392_o = enable_2[130];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4393_o = n4006_o ? 1'b1 : n4392_o;
  assign n4394_o = enable_2[131];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4395_o = n4007_o ? 1'b1 : n4394_o;
  assign n4396_o = enable_2[132];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4397_o = n4008_o ? 1'b1 : n4396_o;
  assign n4398_o = enable_2[133];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4399_o = n4009_o ? 1'b1 : n4398_o;
  assign n4400_o = enable_2[134];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4401_o = n4010_o ? 1'b1 : n4400_o;
  assign n4402_o = enable_2[135];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4403_o = n4011_o ? 1'b1 : n4402_o;
  assign n4404_o = enable_2[136];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4405_o = n4012_o ? 1'b1 : n4404_o;
  assign n4406_o = enable_2[137];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4407_o = n4013_o ? 1'b1 : n4406_o;
  assign n4408_o = enable_2[138];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4409_o = n4014_o ? 1'b1 : n4408_o;
  assign n4410_o = enable_2[139];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4411_o = n4015_o ? 1'b1 : n4410_o;
  assign n4412_o = enable_2[140];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4413_o = n4016_o ? 1'b1 : n4412_o;
  assign n4414_o = enable_2[141];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4415_o = n4017_o ? 1'b1 : n4414_o;
  assign n4416_o = enable_2[142];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4417_o = n4018_o ? 1'b1 : n4416_o;
  assign n4418_o = enable_2[143];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4419_o = n4019_o ? 1'b1 : n4418_o;
  assign n4420_o = enable_2[144];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4421_o = n4020_o ? 1'b1 : n4420_o;
  assign n4422_o = enable_2[145];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4423_o = n4021_o ? 1'b1 : n4422_o;
  assign n4424_o = enable_2[146];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4425_o = n4022_o ? 1'b1 : n4424_o;
  assign n4426_o = enable_2[147];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4427_o = n4023_o ? 1'b1 : n4426_o;
  assign n4428_o = enable_2[148];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4429_o = n4024_o ? 1'b1 : n4428_o;
  assign n4430_o = enable_2[149];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4431_o = n4025_o ? 1'b1 : n4430_o;
  assign n4432_o = enable_2[150];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4433_o = n4026_o ? 1'b1 : n4432_o;
  assign n4434_o = enable_2[151];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4435_o = n4027_o ? 1'b1 : n4434_o;
  assign n4436_o = enable_2[152];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4437_o = n4028_o ? 1'b1 : n4436_o;
  assign n4438_o = enable_2[153];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4439_o = n4029_o ? 1'b1 : n4438_o;
  assign n4440_o = enable_2[154];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4441_o = n4030_o ? 1'b1 : n4440_o;
  assign n4442_o = enable_2[155];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4443_o = n4031_o ? 1'b1 : n4442_o;
  assign n4444_o = enable_2[156];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4445_o = n4032_o ? 1'b1 : n4444_o;
  assign n4446_o = enable_2[157];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4447_o = n4033_o ? 1'b1 : n4446_o;
  assign n4448_o = enable_2[158];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4449_o = n4034_o ? 1'b1 : n4448_o;
  assign n4450_o = enable_2[159];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4451_o = n4035_o ? 1'b1 : n4450_o;
  assign n4452_o = enable_2[160];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4453_o = n4036_o ? 1'b1 : n4452_o;
  assign n4454_o = enable_2[161];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4455_o = n4037_o ? 1'b1 : n4454_o;
  assign n4456_o = enable_2[162];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4457_o = n4038_o ? 1'b1 : n4456_o;
  assign n4458_o = enable_2[163];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4459_o = n4039_o ? 1'b1 : n4458_o;
  assign n4460_o = enable_2[164];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4461_o = n4040_o ? 1'b1 : n4460_o;
  assign n4462_o = enable_2[165];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4463_o = n4041_o ? 1'b1 : n4462_o;
  assign n4464_o = enable_2[166];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4465_o = n4042_o ? 1'b1 : n4464_o;
  assign n4466_o = enable_2[167];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4467_o = n4043_o ? 1'b1 : n4466_o;
  assign n4468_o = enable_2[168];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4469_o = n4044_o ? 1'b1 : n4468_o;
  assign n4470_o = enable_2[169];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4471_o = n4045_o ? 1'b1 : n4470_o;
  assign n4472_o = enable_2[170];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4473_o = n4046_o ? 1'b1 : n4472_o;
  assign n4474_o = enable_2[171];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4475_o = n4047_o ? 1'b1 : n4474_o;
  assign n4476_o = enable_2[172];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4477_o = n4048_o ? 1'b1 : n4476_o;
  assign n4478_o = enable_2[173];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4479_o = n4049_o ? 1'b1 : n4478_o;
  assign n4480_o = enable_2[174];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4481_o = n4050_o ? 1'b1 : n4480_o;
  assign n4482_o = enable_2[175];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4483_o = n4051_o ? 1'b1 : n4482_o;
  assign n4484_o = enable_2[176];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4485_o = n4052_o ? 1'b1 : n4484_o;
  assign n4486_o = enable_2[177];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4487_o = n4053_o ? 1'b1 : n4486_o;
  assign n4488_o = enable_2[178];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4489_o = n4054_o ? 1'b1 : n4488_o;
  assign n4490_o = enable_2[179];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4491_o = n4055_o ? 1'b1 : n4490_o;
  assign n4492_o = enable_2[180];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4493_o = n4056_o ? 1'b1 : n4492_o;
  assign n4494_o = enable_2[181];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4495_o = n4057_o ? 1'b1 : n4494_o;
  assign n4496_o = enable_2[182];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4497_o = n4058_o ? 1'b1 : n4496_o;
  assign n4498_o = enable_2[183];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4499_o = n4059_o ? 1'b1 : n4498_o;
  assign n4500_o = enable_2[184];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4501_o = n4060_o ? 1'b1 : n4500_o;
  assign n4502_o = enable_2[185];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4503_o = n4061_o ? 1'b1 : n4502_o;
  assign n4504_o = enable_2[186];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4505_o = n4062_o ? 1'b1 : n4504_o;
  assign n4506_o = enable_2[187];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4507_o = n4063_o ? 1'b1 : n4506_o;
  assign n4508_o = enable_2[188];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4509_o = n4064_o ? 1'b1 : n4508_o;
  assign n4510_o = enable_2[189];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4511_o = n4065_o ? 1'b1 : n4510_o;
  assign n4512_o = enable_2[190];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4513_o = n4066_o ? 1'b1 : n4512_o;
  assign n4514_o = enable_2[191];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4515_o = n4067_o ? 1'b1 : n4514_o;
  assign n4516_o = enable_2[192];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4517_o = n4068_o ? 1'b1 : n4516_o;
  assign n4518_o = enable_2[193];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4519_o = n4069_o ? 1'b1 : n4518_o;
  assign n4520_o = enable_2[194];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4521_o = n4070_o ? 1'b1 : n4520_o;
  assign n4522_o = enable_2[195];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4523_o = n4071_o ? 1'b1 : n4522_o;
  assign n4524_o = enable_2[196];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4525_o = n4072_o ? 1'b1 : n4524_o;
  assign n4526_o = enable_2[197];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4527_o = n4073_o ? 1'b1 : n4526_o;
  assign n4528_o = enable_2[198];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4529_o = n4074_o ? 1'b1 : n4528_o;
  assign n4530_o = enable_2[199];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4531_o = n4075_o ? 1'b1 : n4530_o;
  assign n4532_o = enable_2[200];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4533_o = n4076_o ? 1'b1 : n4532_o;
  assign n4534_o = enable_2[201];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4535_o = n4077_o ? 1'b1 : n4534_o;
  assign n4536_o = enable_2[202];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4537_o = n4078_o ? 1'b1 : n4536_o;
  assign n4538_o = enable_2[203];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4539_o = n4079_o ? 1'b1 : n4538_o;
  assign n4540_o = enable_2[204];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4541_o = n4080_o ? 1'b1 : n4540_o;
  assign n4542_o = enable_2[205];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4543_o = n4081_o ? 1'b1 : n4542_o;
  assign n4544_o = enable_2[206];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4545_o = n4082_o ? 1'b1 : n4544_o;
  assign n4546_o = enable_2[207];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4547_o = n4083_o ? 1'b1 : n4546_o;
  assign n4548_o = enable_2[208];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4549_o = n4084_o ? 1'b1 : n4548_o;
  assign n4550_o = enable_2[209];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4551_o = n4085_o ? 1'b1 : n4550_o;
  assign n4552_o = enable_2[210];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4553_o = n4086_o ? 1'b1 : n4552_o;
  assign n4554_o = enable_2[211];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4555_o = n4087_o ? 1'b1 : n4554_o;
  assign n4556_o = enable_2[212];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4557_o = n4088_o ? 1'b1 : n4556_o;
  assign n4558_o = enable_2[213];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4559_o = n4089_o ? 1'b1 : n4558_o;
  assign n4560_o = enable_2[214];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4561_o = n4090_o ? 1'b1 : n4560_o;
  assign n4562_o = enable_2[215];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4563_o = n4091_o ? 1'b1 : n4562_o;
  assign n4564_o = enable_2[216];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4565_o = n4092_o ? 1'b1 : n4564_o;
  assign n4566_o = enable_2[217];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4567_o = n4093_o ? 1'b1 : n4566_o;
  assign n4568_o = enable_2[218];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4569_o = n4094_o ? 1'b1 : n4568_o;
  assign n4570_o = enable_2[219];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4571_o = n4095_o ? 1'b1 : n4570_o;
  assign n4572_o = enable_2[220];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4573_o = n4096_o ? 1'b1 : n4572_o;
  assign n4574_o = enable_2[221];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4575_o = n4097_o ? 1'b1 : n4574_o;
  assign n4576_o = enable_2[222];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4577_o = n4098_o ? 1'b1 : n4576_o;
  assign n4578_o = enable_2[223];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4579_o = n4099_o ? 1'b1 : n4578_o;
  assign n4580_o = enable_2[224];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4581_o = n4100_o ? 1'b1 : n4580_o;
  assign n4582_o = enable_2[225];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4583_o = n4101_o ? 1'b1 : n4582_o;
  assign n4584_o = enable_2[226];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4585_o = n4102_o ? 1'b1 : n4584_o;
  assign n4586_o = enable_2[227];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4587_o = n4103_o ? 1'b1 : n4586_o;
  assign n4588_o = enable_2[228];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4589_o = n4104_o ? 1'b1 : n4588_o;
  assign n4590_o = enable_2[229];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4591_o = n4105_o ? 1'b1 : n4590_o;
  assign n4592_o = enable_2[230];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4593_o = n4106_o ? 1'b1 : n4592_o;
  assign n4594_o = enable_2[231];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4595_o = n4107_o ? 1'b1 : n4594_o;
  assign n4596_o = enable_2[232];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4597_o = n4108_o ? 1'b1 : n4596_o;
  assign n4598_o = enable_2[233];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4599_o = n4109_o ? 1'b1 : n4598_o;
  assign n4600_o = enable_2[234];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4601_o = n4110_o ? 1'b1 : n4600_o;
  assign n4602_o = enable_2[235];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4603_o = n4111_o ? 1'b1 : n4602_o;
  assign n4604_o = enable_2[236];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4605_o = n4112_o ? 1'b1 : n4604_o;
  assign n4606_o = enable_2[237];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4607_o = n4113_o ? 1'b1 : n4606_o;
  assign n4608_o = enable_2[238];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4609_o = n4114_o ? 1'b1 : n4608_o;
  assign n4610_o = enable_2[239];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4611_o = n4115_o ? 1'b1 : n4610_o;
  assign n4612_o = enable_2[240];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4613_o = n4116_o ? 1'b1 : n4612_o;
  assign n4614_o = enable_2[241];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4615_o = n4117_o ? 1'b1 : n4614_o;
  assign n4616_o = enable_2[242];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4617_o = n4118_o ? 1'b1 : n4616_o;
  assign n4618_o = enable_2[243];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4619_o = n4119_o ? 1'b1 : n4618_o;
  assign n4620_o = enable_2[244];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4621_o = n4120_o ? 1'b1 : n4620_o;
  assign n4622_o = enable_2[245];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4623_o = n4121_o ? 1'b1 : n4622_o;
  assign n4624_o = enable_2[246];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4625_o = n4122_o ? 1'b1 : n4624_o;
  assign n4626_o = enable_2[247];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4627_o = n4123_o ? 1'b1 : n4626_o;
  assign n4628_o = enable_2[248];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4629_o = n4124_o ? 1'b1 : n4628_o;
  assign n4630_o = enable_2[249];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4631_o = n4125_o ? 1'b1 : n4630_o;
  assign n4632_o = enable_2[250];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4633_o = n4126_o ? 1'b1 : n4632_o;
  assign n4634_o = enable_2[251];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4635_o = n4127_o ? 1'b1 : n4634_o;
  assign n4636_o = enable_2[252];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4637_o = n4128_o ? 1'b1 : n4636_o;
  assign n4638_o = enable_2[253];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4639_o = n4129_o ? 1'b1 : n4638_o;
  assign n4640_o = enable_2[254];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4641_o = n4130_o ? 1'b1 : n4640_o;
  assign n4642_o = enable_2[255];
  /* RTL_PUF/vhdl/ro_puf_s7.vhd:438:21  */
  assign n4643_o = n4131_o ? 1'b1 : n4642_o;
  assign n4644_o = {n4643_o, n4641_o, n4639_o, n4637_o, n4635_o, n4633_o, n4631_o, n4629_o, n4627_o, n4625_o, n4623_o, n4621_o, n4619_o, n4617_o, n4615_o, n4613_o, n4611_o, n4609_o, n4607_o, n4605_o, n4603_o, n4601_o, n4599_o, n4597_o, n4595_o, n4593_o, n4591_o, n4589_o, n4587_o, n4585_o, n4583_o, n4581_o, n4579_o, n4577_o, n4575_o, n4573_o, n4571_o, n4569_o, n4567_o, n4565_o, n4563_o, n4561_o, n4559_o, n4557_o, n4555_o, n4553_o, n4551_o, n4549_o, n4547_o, n4545_o, n4543_o, n4541_o, n4539_o, n4537_o, n4535_o, n4533_o, n4531_o, n4529_o, n4527_o, n4525_o, n4523_o, n4521_o, n4519_o, n4517_o, n4515_o, n4513_o, n4511_o, n4509_o, n4507_o, n4505_o, n4503_o, n4501_o, n4499_o, n4497_o, n4495_o, n4493_o, n4491_o, n4489_o, n4487_o, n4485_o, n4483_o, n4481_o, n4479_o, n4477_o, n4475_o, n4473_o, n4471_o, n4469_o, n4467_o, n4465_o, n4463_o, n4461_o, n4459_o, n4457_o, n4455_o, n4453_o, n4451_o, n4449_o, n4447_o, n4445_o, n4443_o, n4441_o, n4439_o, n4437_o, n4435_o, n4433_o, n4431_o, n4429_o, n4427_o, n4425_o, n4423_o, n4421_o, n4419_o, n4417_o, n4415_o, n4413_o, n4411_o, n4409_o, n4407_o, n4405_o, n4403_o, n4401_o, n4399_o, n4397_o, n4395_o, n4393_o, n4391_o, n4389_o, n4387_o, n4385_o, n4383_o, n4381_o, n4379_o, n4377_o, n4375_o, n4373_o, n4371_o, n4369_o, n4367_o, n4365_o, n4363_o, n4361_o, n4359_o, n4357_o, n4355_o, n4353_o, n4351_o, n4349_o, n4347_o, n4345_o, n4343_o, n4341_o, n4339_o, n4337_o, n4335_o, n4333_o, n4331_o, n4329_o, n4327_o, n4325_o, n4323_o, n4321_o, n4319_o, n4317_o, n4315_o, n4313_o, n4311_o, n4309_o, n4307_o, n4305_o, n4303_o, n4301_o, n4299_o, n4297_o, n4295_o, n4293_o, n4291_o, n4289_o, n4287_o, n4285_o, n4283_o, n4281_o, n4279_o, n4277_o, n4275_o, n4273_o, n4271_o, n4269_o, n4267_o, n4265_o, n4263_o, n4261_o, n4259_o, n4257_o, n4255_o, n4253_o, n4251_o, n4249_o, n4247_o, n4245_o, n4243_o, n4241_o, n4239_o, n4237_o, n4235_o, n4233_o, n4231_o, n4229_o, n4227_o, n4225_o, n4223_o, n4221_o, n4219_o, n4217_o, n4215_o, n4213_o, n4211_o, n4209_o, n4207_o, n4205_o, n4203_o, n4201_o, n4199_o, n4197_o, n4195_o, n4193_o, n4191_o, n4189_o, n4187_o, n4185_o, n4183_o, n4181_o, n4179_o, n4177_o, n4175_o, n4173_o, n4171_o, n4169_o, n4167_o, n4165_o, n4163_o, n4161_o, n4159_o, n4157_o, n4155_o, n4153_o, n4151_o, n4149_o, n4147_o, n4145_o, n4143_o, n4141_o, n4139_o, n4137_o, n4135_o, n4133_o};
endmodule

